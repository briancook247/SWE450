// Computer_System.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module Computer_System (
		output wire        adc_sclk,                        //                  adc.sclk
		output wire        adc_cs_n,                        //                     .cs_n
		input  wire        adc_dout,                        //                     .dout
		output wire        adc_din,                         //                     .din
		input  wire        audio_ADCDAT,                    //                audio.ADCDAT
		input  wire        audio_ADCLRCK,                   //                     .ADCLRCK
		input  wire        audio_BCLK,                      //                     .BCLK
		output wire        audio_DACDAT,                    //                     .DACDAT
		input  wire        audio_DACLRCK,                   //                     .DACLRCK
		output wire        audio_pll_clk_clk,               //        audio_pll_clk.clk
		input  wire        audio_pll_ref_clk_clk,           //    audio_pll_ref_clk.clk
		input  wire        audio_pll_ref_reset_reset,       //  audio_pll_ref_reset.reset
		inout  wire        av_config_SDAT,                  //            av_config.SDAT
		output wire        av_config_SCLK,                  //                     .SCLK
		inout  wire [31:0] expansion_jp1_export,            //        expansion_jp1.export
		output wire [31:0] hex3_hex0_export,                //            hex3_hex0.export
		output wire [15:0] hex5_hex4_export,                //            hex5_hex4.export
		output wire        hps_io_hps_io_emac1_inst_TX_CLK, //               hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,   //                     .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,   //                     .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,   //                     .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,   //                     .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,   //                     .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,   //                     .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,    //                     .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL, //                     .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL, //                     .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK, //                     .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,   //                     .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,   //                     .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,   //                     .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_qspi_inst_IO0,     //                     .hps_io_qspi_inst_IO0
		inout  wire        hps_io_hps_io_qspi_inst_IO1,     //                     .hps_io_qspi_inst_IO1
		inout  wire        hps_io_hps_io_qspi_inst_IO2,     //                     .hps_io_qspi_inst_IO2
		inout  wire        hps_io_hps_io_qspi_inst_IO3,     //                     .hps_io_qspi_inst_IO3
		output wire        hps_io_hps_io_qspi_inst_SS0,     //                     .hps_io_qspi_inst_SS0
		output wire        hps_io_hps_io_qspi_inst_CLK,     //                     .hps_io_qspi_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_CMD,     //                     .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,      //                     .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,      //                     .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,     //                     .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,      //                     .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,      //                     .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,      //                     .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,      //                     .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,      //                     .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,      //                     .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,      //                     .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,      //                     .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,      //                     .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,      //                     .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,     //                     .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,     //                     .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,     //                     .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,     //                     .hps_io_usb1_inst_NXT
		output wire        hps_io_hps_io_spim0_inst_CLK,    //                     .hps_io_spim0_inst_CLK
		output wire        hps_io_hps_io_spim0_inst_MOSI,   //                     .hps_io_spim0_inst_MOSI
		input  wire        hps_io_hps_io_spim0_inst_MISO,   //                     .hps_io_spim0_inst_MISO
		output wire        hps_io_hps_io_spim0_inst_SS0,    //                     .hps_io_spim0_inst_SS0
		output wire        hps_io_hps_io_spim1_inst_CLK,    //                     .hps_io_spim1_inst_CLK
		output wire        hps_io_hps_io_spim1_inst_MOSI,   //                     .hps_io_spim1_inst_MOSI
		input  wire        hps_io_hps_io_spim1_inst_MISO,   //                     .hps_io_spim1_inst_MISO
		output wire        hps_io_hps_io_spim1_inst_SS0,    //                     .hps_io_spim1_inst_SS0
		input  wire        hps_io_hps_io_uart0_inst_RX,     //                     .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,     //                     .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,     //                     .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,     //                     .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,     //                     .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,     //                     .hps_io_i2c1_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,  //                     .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,  //                     .hps_io_gpio_inst_GPIO35
		inout  wire        hps_io_hps_io_gpio_inst_GPIO37,  //                     .hps_io_gpio_inst_GPIO37
		inout  wire        hps_io_hps_io_gpio_inst_GPIO40,  //                     .hps_io_gpio_inst_GPIO40
		inout  wire        hps_io_hps_io_gpio_inst_GPIO41,  //                     .hps_io_gpio_inst_GPIO41
		inout  wire        hps_io_hps_io_gpio_inst_GPIO44,  //                     .hps_io_gpio_inst_GPIO44
		inout  wire        hps_io_hps_io_gpio_inst_GPIO48,  //                     .hps_io_gpio_inst_GPIO48
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53,  //                     .hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54,  //                     .hps_io_gpio_inst_GPIO54
		inout  wire        hps_io_hps_io_gpio_inst_GPIO61,  //                     .hps_io_gpio_inst_GPIO61
		output wire        irda_TXD,                        //                 irda.TXD
		input  wire        irda_RXD,                        //                     .RXD
		output wire [9:0]  leds_export,                     //                 leds.export
		output wire [14:0] memory_mem_a,                    //               memory.mem_a
		output wire [2:0]  memory_mem_ba,                   //                     .mem_ba
		output wire        memory_mem_ck,                   //                     .mem_ck
		output wire        memory_mem_ck_n,                 //                     .mem_ck_n
		output wire        memory_mem_cke,                  //                     .mem_cke
		output wire        memory_mem_cs_n,                 //                     .mem_cs_n
		output wire        memory_mem_ras_n,                //                     .mem_ras_n
		output wire        memory_mem_cas_n,                //                     .mem_cas_n
		output wire        memory_mem_we_n,                 //                     .mem_we_n
		output wire        memory_mem_reset_n,              //                     .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                   //                     .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                  //                     .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                //                     .mem_dqs_n
		output wire        memory_mem_odt,                  //                     .mem_odt
		output wire [3:0]  memory_mem_dm,                   //                     .mem_dm
		input  wire        memory_oct_rzqin,                //                     .oct_rzqin
		inout  wire        ps2_port_CLK,                    //             ps2_port.CLK
		inout  wire        ps2_port_DAT,                    //                     .DAT
		inout  wire        ps2_port_dual_CLK,               //        ps2_port_dual.CLK
		inout  wire        ps2_port_dual_DAT,               //                     .DAT
		input  wire [3:0]  pushbuttons_export,              //          pushbuttons.export
		output wire [12:0] sdram_addr,                      //                sdram.addr
		output wire [1:0]  sdram_ba,                        //                     .ba
		output wire        sdram_cas_n,                     //                     .cas_n
		output wire        sdram_cke,                       //                     .cke
		output wire        sdram_cs_n,                      //                     .cs_n
		inout  wire [15:0] sdram_dq,                        //                     .dq
		output wire [1:0]  sdram_dqm,                       //                     .dqm
		output wire        sdram_ras_n,                     //                     .ras_n
		output wire        sdram_we_n,                      //                     .we_n
		output wire        sdram_clk_clk,                   //            sdram_clk.clk
		input  wire [9:0]  slider_switches_export,          //      slider_switches.export
		input  wire        system_pll_ref_clk_clk,          //   system_pll_ref_clk.clk
		input  wire        system_pll_ref_reset_reset,      // system_pll_ref_reset.reset
		output wire        vga_CLK,                         //                  vga.CLK
		output wire        vga_HS,                          //                     .HS
		output wire        vga_VS,                          //                     .VS
		output wire        vga_BLANK,                       //                     .BLANK
		output wire        vga_SYNC,                        //                     .SYNC
		output wire [7:0]  vga_R,                           //                     .R
		output wire [7:0]  vga_G,                           //                     .G
		output wire [7:0]  vga_B,                           //                     .B
		input  wire        video_in_TD_CLK27,               //             video_in.TD_CLK27
		input  wire [7:0]  video_in_TD_DATA,                //                     .TD_DATA
		input  wire        video_in_TD_HS,                  //                     .TD_HS
		input  wire        video_in_TD_VS,                  //                     .TD_VS
		input  wire        video_in_clk27_reset,            //                     .clk27_reset
		output wire        video_in_TD_RESET,               //                     .TD_RESET
		output wire        video_in_overflow_flag,          //                     .overflow_flag
		input  wire        video_pll_ref_clk_clk,           //    video_pll_ref_clk.clk
		input  wire        video_pll_ref_reset_reset        //  video_pll_ref_reset.reset
	);

	wire         system_pll_sys_clk_clk;                                                                // System_PLL:sys_clk_clk -> [ADC:clock, ARM_A9_HPS:f2h_axi_clk, ARM_A9_HPS:h2f_axi_clk, ARM_A9_HPS:h2f_lw_axi_clk, AV_Config:clk, Audio_Subsystem:sys_clk_clk, Char_DMA_Addr_Translation:clk, Expansion_JP1:clk, F2H_Mem_Window_00000000:clk, F2H_Mem_Window_FF600000:clk, F2H_Mem_Window_FF800000:clk, HEX3_HEX0:clk, HEX5_HEX4:clk, Interval_Timer:clk, Interval_Timer_2:clk, Interval_Timer_2nd_Core:clk, Interval_Timer_2nd_Core_2:clk, IrDA:clk, JTAG_UART:clk, JTAG_UART_2nd_Core:clk, JTAG_UART_for_ARM_0:clk, JTAG_UART_for_ARM_1:clk, JTAG_to_FPGA_Bridge:clk_clk, JTAG_to_HPS_Bridge:clk_clk, LEDs:clk, Nios2:clk, Nios2_2nd_Core:clk, Onchip_SRAM:clk, PS2_Port:clk, PS2_Port_Dual:clk, Pixel_DMA_Addr_Translation:clk, Pushbuttons:clk, SDRAM:clk, Slider_Switches:clk, SysID:clock, VGA_Subsystem:sys_clk_clk, Video_In_DMA_Addr_Translation:clk, Video_In_Subsystem:sys_clk_clk, irq_mapper_002:clk, irq_mapper_003:clk, mm_interconnect_0:System_PLL_sys_clk_clk, mm_interconnect_1:System_PLL_sys_clk_clk, rst_controller:clk, rst_controller_004:clk, rst_controller_005:clk, rst_controller_008:clk]
	wire         video_pll_vga_clk_clk;                                                                 // Video_PLL:vga_clk_clk -> VGA_Subsystem:vga_clk_clk
	wire         video_pll_reset_source_reset;                                                          // Video_PLL:reset_source_reset -> VGA_Subsystem:vga_reset_reset_n
	wire  [31:0] nios2_custom_instruction_master_multi_dataa;                                           // Nios2:A_ci_multi_dataa -> Nios2_custom_instruction_master_translator:ci_slave_multi_dataa
	wire         nios2_custom_instruction_master_multi_writerc;                                         // Nios2:A_ci_multi_writerc -> Nios2_custom_instruction_master_translator:ci_slave_multi_writerc
	wire  [31:0] nios2_custom_instruction_master_multi_result;                                          // Nios2_custom_instruction_master_translator:ci_slave_multi_result -> Nios2:A_ci_multi_result
	wire         nios2_custom_instruction_master_clk;                                                   // Nios2:A_ci_multi_clock -> Nios2_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] nios2_custom_instruction_master_multi_datab;                                           // Nios2:A_ci_multi_datab -> Nios2_custom_instruction_master_translator:ci_slave_multi_datab
	wire         nios2_custom_instruction_master_start;                                                 // Nios2:A_ci_multi_start -> Nios2_custom_instruction_master_translator:ci_slave_multi_start
	wire   [4:0] nios2_custom_instruction_master_multi_b;                                               // Nios2:A_ci_multi_b -> Nios2_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] nios2_custom_instruction_master_multi_c;                                               // Nios2:A_ci_multi_c -> Nios2_custom_instruction_master_translator:ci_slave_multi_c
	wire         nios2_custom_instruction_master_reset_req;                                             // Nios2:A_ci_multi_reset_req -> Nios2_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         nios2_custom_instruction_master_done;                                                  // Nios2_custom_instruction_master_translator:ci_slave_multi_done -> Nios2:A_ci_multi_done
	wire   [4:0] nios2_custom_instruction_master_multi_a;                                               // Nios2:A_ci_multi_a -> Nios2_custom_instruction_master_translator:ci_slave_multi_a
	wire         nios2_custom_instruction_master_clk_en;                                                // Nios2:A_ci_multi_clk_en -> Nios2_custom_instruction_master_translator:ci_slave_multi_clken
	wire         nios2_custom_instruction_master_reset;                                                 // Nios2:A_ci_multi_reset -> Nios2_custom_instruction_master_translator:ci_slave_multi_reset
	wire         nios2_custom_instruction_master_multi_readrb;                                          // Nios2:A_ci_multi_readrb -> Nios2_custom_instruction_master_translator:ci_slave_multi_readrb
	wire         nios2_custom_instruction_master_multi_readra;                                          // Nios2:A_ci_multi_readra -> Nios2_custom_instruction_master_translator:ci_slave_multi_readra
	wire   [7:0] nios2_custom_instruction_master_multi_n;                                               // Nios2:A_ci_multi_n -> Nios2_custom_instruction_master_translator:ci_slave_multi_n
	wire         nios2_custom_instruction_master_translator_multi_ci_master_readra;                     // Nios2_custom_instruction_master_translator:multi_ci_master_readra -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] nios2_custom_instruction_master_translator_multi_ci_master_a;                          // Nios2_custom_instruction_master_translator:multi_ci_master_a -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] nios2_custom_instruction_master_translator_multi_ci_master_b;                          // Nios2_custom_instruction_master_translator:multi_ci_master_b -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         nios2_custom_instruction_master_translator_multi_ci_master_clk;                        // Nios2_custom_instruction_master_translator:multi_ci_master_clk -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios2_custom_instruction_master_translator_multi_ci_master_readrb;                     // Nios2_custom_instruction_master_translator:multi_ci_master_readrb -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] nios2_custom_instruction_master_translator_multi_ci_master_c;                          // Nios2_custom_instruction_master_translator:multi_ci_master_c -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         nios2_custom_instruction_master_translator_multi_ci_master_start;                      // Nios2_custom_instruction_master_translator:multi_ci_master_start -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         nios2_custom_instruction_master_translator_multi_ci_master_reset_req;                  // Nios2_custom_instruction_master_translator:multi_ci_master_reset_req -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios2_custom_instruction_master_translator_multi_ci_master_done;                       // Nios2_custom_instruction_master_multi_xconnect:ci_slave_done -> Nios2_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios2_custom_instruction_master_translator_multi_ci_master_n;                          // Nios2_custom_instruction_master_translator:multi_ci_master_n -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] nios2_custom_instruction_master_translator_multi_ci_master_result;                     // Nios2_custom_instruction_master_multi_xconnect:ci_slave_result -> Nios2_custom_instruction_master_translator:multi_ci_master_result
	wire         nios2_custom_instruction_master_translator_multi_ci_master_clk_en;                     // Nios2_custom_instruction_master_translator:multi_ci_master_clken -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] nios2_custom_instruction_master_translator_multi_ci_master_datab;                      // Nios2_custom_instruction_master_translator:multi_ci_master_datab -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] nios2_custom_instruction_master_translator_multi_ci_master_dataa;                      // Nios2_custom_instruction_master_translator:multi_ci_master_dataa -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios2_custom_instruction_master_translator_multi_ci_master_reset;                      // Nios2_custom_instruction_master_translator:multi_ci_master_reset -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         nios2_custom_instruction_master_translator_multi_ci_master_writerc;                    // Nios2_custom_instruction_master_translator:multi_ci_master_writerc -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_readra;                      // Nios2_custom_instruction_master_multi_xconnect:ci_master0_readra -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_a;                           // Nios2_custom_instruction_master_multi_xconnect:ci_master0_a -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_b;                           // Nios2_custom_instruction_master_multi_xconnect:ci_master0_b -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_readrb;                      // Nios2_custom_instruction_master_multi_xconnect:ci_master0_readrb -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_c;                           // Nios2_custom_instruction_master_multi_xconnect:ci_master0_c -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_clk;                         // Nios2_custom_instruction_master_multi_xconnect:ci_master0_clk -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_ipending;                    // Nios2_custom_instruction_master_multi_xconnect:ci_master0_ipending -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_start;                       // Nios2_custom_instruction_master_multi_xconnect:ci_master0_start -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_reset_req;                   // Nios2_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_done;                        // Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_done -> Nios2_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_n;                           // Nios2_custom_instruction_master_multi_xconnect:ci_master0_n -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_result;                      // Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_result -> Nios2_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_estatus;                     // Nios2_custom_instruction_master_multi_xconnect:ci_master0_estatus -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_clk_en;                      // Nios2_custom_instruction_master_multi_xconnect:ci_master0_clken -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_datab;                       // Nios2_custom_instruction_master_multi_xconnect:ci_master0_datab -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_dataa;                       // Nios2_custom_instruction_master_multi_xconnect:ci_master0_dataa -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_reset;                       // Nios2_custom_instruction_master_multi_xconnect:ci_master0_reset -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_writerc;                     // Nios2_custom_instruction_master_multi_xconnect:ci_master0_writerc -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios2_custom_instruction_master_multi_slave_translator0_ci_master_result;              // Nios2_Floating_Point:result -> Nios2_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk;                 // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_clk -> Nios2_Floating_Point:clk
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;              // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_clken -> Nios2_Floating_Point:clk_en
	wire  [31:0] nios2_custom_instruction_master_multi_slave_translator0_ci_master_datab;               // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_datab -> Nios2_Floating_Point:datab
	wire  [31:0] nios2_custom_instruction_master_multi_slave_translator0_ci_master_dataa;               // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> Nios2_Floating_Point:dataa
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_start;               // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_start -> Nios2_Floating_Point:start
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_reset;               // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_reset -> Nios2_Floating_Point:reset
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_done;                // Nios2_Floating_Point:done -> Nios2_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [1:0] nios2_custom_instruction_master_multi_slave_translator0_ci_master_n;                   // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_n -> Nios2_Floating_Point:n
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_dataa;                                  // Nios2_2nd_Core:A_ci_multi_dataa -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_dataa
	wire         nios2_2nd_core_custom_instruction_master_multi_writerc;                                // Nios2_2nd_Core:A_ci_multi_writerc -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_writerc
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_result;                                 // Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_result -> Nios2_2nd_Core:A_ci_multi_result
	wire         nios2_2nd_core_custom_instruction_master_clk;                                          // Nios2_2nd_Core:A_ci_multi_clock -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_datab;                                  // Nios2_2nd_Core:A_ci_multi_datab -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_datab
	wire         nios2_2nd_core_custom_instruction_master_start;                                        // Nios2_2nd_Core:A_ci_multi_start -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_start
	wire   [4:0] nios2_2nd_core_custom_instruction_master_multi_b;                                      // Nios2_2nd_Core:A_ci_multi_b -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] nios2_2nd_core_custom_instruction_master_multi_c;                                      // Nios2_2nd_Core:A_ci_multi_c -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_c
	wire         nios2_2nd_core_custom_instruction_master_reset_req;                                    // Nios2_2nd_Core:A_ci_multi_reset_req -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         nios2_2nd_core_custom_instruction_master_done;                                         // Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_done -> Nios2_2nd_Core:A_ci_multi_done
	wire   [4:0] nios2_2nd_core_custom_instruction_master_multi_a;                                      // Nios2_2nd_Core:A_ci_multi_a -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_a
	wire         nios2_2nd_core_custom_instruction_master_clk_en;                                       // Nios2_2nd_Core:A_ci_multi_clk_en -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_clken
	wire         nios2_2nd_core_custom_instruction_master_reset;                                        // Nios2_2nd_Core:A_ci_multi_reset -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_reset
	wire         nios2_2nd_core_custom_instruction_master_multi_readrb;                                 // Nios2_2nd_Core:A_ci_multi_readrb -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_readrb
	wire         nios2_2nd_core_custom_instruction_master_multi_readra;                                 // Nios2_2nd_Core:A_ci_multi_readra -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_readra
	wire   [7:0] nios2_2nd_core_custom_instruction_master_multi_n;                                      // Nios2_2nd_Core:A_ci_multi_n -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_n
	wire         nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_readra;            // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_readra -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_a;                 // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_a -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_b;                 // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_b -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_clk;               // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_clk -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_readrb;            // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_readrb -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_c;                 // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_c -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_start;             // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_start -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_reset_req;         // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_reset_req -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_done;              // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_done -> Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_n;                 // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_n -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_result;            // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_result -> Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_result
	wire         nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_clk_en;            // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_clken -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_datab;             // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_datab -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_dataa;             // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_dataa -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_reset;             // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_reset -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_writerc;           // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_writerc -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_readra;             // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_readra -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_a;                  // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_a -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_b;                  // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_b -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_readrb;             // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_readrb -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_c;                  // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_c -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_clk;                // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_clk -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_ipending;           // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_ipending -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_start;              // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_start -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_reset_req;          // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_done;               // Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_done -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_n;                  // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_n -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_result;             // Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_result -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_estatus;            // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_estatus -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_clk_en;             // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_clken -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_datab;              // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_datab -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_dataa;              // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_dataa -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_reset;              // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_reset -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_writerc;            // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_writerc -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_result;     // Nios2_2nd_Core_Floating_Point:result -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_clk;        // Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_master_clk -> Nios2_2nd_Core_Floating_Point:clk
	wire         nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;     // Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_master_clken -> Nios2_2nd_Core_Floating_Point:clk_en
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_datab;      // Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_master_datab -> Nios2_2nd_Core_Floating_Point:datab
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_dataa;      // Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> Nios2_2nd_Core_Floating_Point:dataa
	wire         nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_start;      // Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_master_start -> Nios2_2nd_Core_Floating_Point:start
	wire         nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_reset;      // Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_master_reset -> Nios2_2nd_Core_Floating_Point:reset
	wire         nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_done;       // Nios2_2nd_Core_Floating_Point:done -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [1:0] nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_n;          // Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_master_n -> Nios2_2nd_Core_Floating_Point:n
	wire  [31:0] nios2_data_master_readdata;                                                            // mm_interconnect_0:Nios2_data_master_readdata -> Nios2:d_readdata
	wire         nios2_data_master_waitrequest;                                                         // mm_interconnect_0:Nios2_data_master_waitrequest -> Nios2:d_waitrequest
	wire         nios2_data_master_debugaccess;                                                         // Nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Nios2_data_master_debugaccess
	wire  [31:0] nios2_data_master_address;                                                             // Nios2:d_address -> mm_interconnect_0:Nios2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                                                          // Nios2:d_byteenable -> mm_interconnect_0:Nios2_data_master_byteenable
	wire         nios2_data_master_read;                                                                // Nios2:d_read -> mm_interconnect_0:Nios2_data_master_read
	wire         nios2_data_master_write;                                                               // Nios2:d_write -> mm_interconnect_0:Nios2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                                                           // Nios2:d_writedata -> mm_interconnect_0:Nios2_data_master_writedata
	wire  [31:0] nios2_2nd_core_data_master_readdata;                                                   // mm_interconnect_0:Nios2_2nd_Core_data_master_readdata -> Nios2_2nd_Core:d_readdata
	wire         nios2_2nd_core_data_master_waitrequest;                                                // mm_interconnect_0:Nios2_2nd_Core_data_master_waitrequest -> Nios2_2nd_Core:d_waitrequest
	wire         nios2_2nd_core_data_master_debugaccess;                                                // Nios2_2nd_Core:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Nios2_2nd_Core_data_master_debugaccess
	wire  [31:0] nios2_2nd_core_data_master_address;                                                    // Nios2_2nd_Core:d_address -> mm_interconnect_0:Nios2_2nd_Core_data_master_address
	wire   [3:0] nios2_2nd_core_data_master_byteenable;                                                 // Nios2_2nd_Core:d_byteenable -> mm_interconnect_0:Nios2_2nd_Core_data_master_byteenable
	wire         nios2_2nd_core_data_master_read;                                                       // Nios2_2nd_Core:d_read -> mm_interconnect_0:Nios2_2nd_Core_data_master_read
	wire         nios2_2nd_core_data_master_write;                                                      // Nios2_2nd_Core:d_write -> mm_interconnect_0:Nios2_2nd_Core_data_master_write
	wire  [31:0] nios2_2nd_core_data_master_writedata;                                                  // Nios2_2nd_Core:d_writedata -> mm_interconnect_0:Nios2_2nd_Core_data_master_writedata
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_awburst;                                                  // ARM_A9_HPS:h2f_lw_AWBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awburst
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_arlen;                                                    // ARM_A9_HPS:h2f_lw_ARLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arlen
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_wstrb;                                                    // ARM_A9_HPS:h2f_lw_WSTRB -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wstrb
	wire         arm_a9_hps_h2f_lw_axi_master_wready;                                                   // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wready -> ARM_A9_HPS:h2f_lw_WREADY
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_rid;                                                      // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rid -> ARM_A9_HPS:h2f_lw_RID
	wire         arm_a9_hps_h2f_lw_axi_master_rready;                                                   // ARM_A9_HPS:h2f_lw_RREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rready
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_awlen;                                                    // ARM_A9_HPS:h2f_lw_AWLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awlen
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_wid;                                                      // ARM_A9_HPS:h2f_lw_WID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wid
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_arcache;                                                  // ARM_A9_HPS:h2f_lw_ARCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arcache
	wire         arm_a9_hps_h2f_lw_axi_master_wvalid;                                                   // ARM_A9_HPS:h2f_lw_WVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wvalid
	wire  [20:0] arm_a9_hps_h2f_lw_axi_master_araddr;                                                   // ARM_A9_HPS:h2f_lw_ARADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_araddr
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_arprot;                                                   // ARM_A9_HPS:h2f_lw_ARPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arprot
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_awprot;                                                   // ARM_A9_HPS:h2f_lw_AWPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awprot
	wire  [31:0] arm_a9_hps_h2f_lw_axi_master_wdata;                                                    // ARM_A9_HPS:h2f_lw_WDATA -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wdata
	wire         arm_a9_hps_h2f_lw_axi_master_arvalid;                                                  // ARM_A9_HPS:h2f_lw_ARVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arvalid
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_awcache;                                                  // ARM_A9_HPS:h2f_lw_AWCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awcache
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_arid;                                                     // ARM_A9_HPS:h2f_lw_ARID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arid
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_arlock;                                                   // ARM_A9_HPS:h2f_lw_ARLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arlock
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_awlock;                                                   // ARM_A9_HPS:h2f_lw_AWLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awlock
	wire  [20:0] arm_a9_hps_h2f_lw_axi_master_awaddr;                                                   // ARM_A9_HPS:h2f_lw_AWADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awaddr
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_bresp;                                                    // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bresp -> ARM_A9_HPS:h2f_lw_BRESP
	wire         arm_a9_hps_h2f_lw_axi_master_arready;                                                  // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arready -> ARM_A9_HPS:h2f_lw_ARREADY
	wire  [31:0] arm_a9_hps_h2f_lw_axi_master_rdata;                                                    // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rdata -> ARM_A9_HPS:h2f_lw_RDATA
	wire         arm_a9_hps_h2f_lw_axi_master_awready;                                                  // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awready -> ARM_A9_HPS:h2f_lw_AWREADY
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_arburst;                                                  // ARM_A9_HPS:h2f_lw_ARBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arburst
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_arsize;                                                   // ARM_A9_HPS:h2f_lw_ARSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arsize
	wire         arm_a9_hps_h2f_lw_axi_master_bready;                                                   // ARM_A9_HPS:h2f_lw_BREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bready
	wire         arm_a9_hps_h2f_lw_axi_master_rlast;                                                    // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rlast -> ARM_A9_HPS:h2f_lw_RLAST
	wire         arm_a9_hps_h2f_lw_axi_master_wlast;                                                    // ARM_A9_HPS:h2f_lw_WLAST -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wlast
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_rresp;                                                    // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rresp -> ARM_A9_HPS:h2f_lw_RRESP
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_awid;                                                     // ARM_A9_HPS:h2f_lw_AWID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awid
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_bid;                                                      // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bid -> ARM_A9_HPS:h2f_lw_BID
	wire         arm_a9_hps_h2f_lw_axi_master_bvalid;                                                   // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bvalid -> ARM_A9_HPS:h2f_lw_BVALID
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_awsize;                                                   // ARM_A9_HPS:h2f_lw_AWSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awsize
	wire         arm_a9_hps_h2f_lw_axi_master_awvalid;                                                  // ARM_A9_HPS:h2f_lw_AWVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awvalid
	wire         arm_a9_hps_h2f_lw_axi_master_rvalid;                                                   // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rvalid -> ARM_A9_HPS:h2f_lw_RVALID
	wire  [31:0] jtag_to_fpga_bridge_master_readdata;                                                   // mm_interconnect_0:JTAG_to_FPGA_Bridge_master_readdata -> JTAG_to_FPGA_Bridge:master_readdata
	wire         jtag_to_fpga_bridge_master_waitrequest;                                                // mm_interconnect_0:JTAG_to_FPGA_Bridge_master_waitrequest -> JTAG_to_FPGA_Bridge:master_waitrequest
	wire  [31:0] jtag_to_fpga_bridge_master_address;                                                    // JTAG_to_FPGA_Bridge:master_address -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_address
	wire         jtag_to_fpga_bridge_master_read;                                                       // JTAG_to_FPGA_Bridge:master_read -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_read
	wire   [3:0] jtag_to_fpga_bridge_master_byteenable;                                                 // JTAG_to_FPGA_Bridge:master_byteenable -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_byteenable
	wire         jtag_to_fpga_bridge_master_readdatavalid;                                              // mm_interconnect_0:JTAG_to_FPGA_Bridge_master_readdatavalid -> JTAG_to_FPGA_Bridge:master_readdatavalid
	wire         jtag_to_fpga_bridge_master_write;                                                      // JTAG_to_FPGA_Bridge:master_write -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_write
	wire  [31:0] jtag_to_fpga_bridge_master_writedata;                                                  // JTAG_to_FPGA_Bridge:master_writedata -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_writedata
	wire  [31:0] video_in_dma_addr_translation_master_readdata;                                         // mm_interconnect_0:Video_In_DMA_Addr_Translation_master_readdata -> Video_In_DMA_Addr_Translation:master_readdata
	wire         video_in_dma_addr_translation_master_waitrequest;                                      // mm_interconnect_0:Video_In_DMA_Addr_Translation_master_waitrequest -> Video_In_DMA_Addr_Translation:master_waitrequest
	wire   [1:0] video_in_dma_addr_translation_master_address;                                          // Video_In_DMA_Addr_Translation:master_address -> mm_interconnect_0:Video_In_DMA_Addr_Translation_master_address
	wire   [3:0] video_in_dma_addr_translation_master_byteenable;                                       // Video_In_DMA_Addr_Translation:master_byteenable -> mm_interconnect_0:Video_In_DMA_Addr_Translation_master_byteenable
	wire         video_in_dma_addr_translation_master_read;                                             // Video_In_DMA_Addr_Translation:master_read -> mm_interconnect_0:Video_In_DMA_Addr_Translation_master_read
	wire         video_in_dma_addr_translation_master_write;                                            // Video_In_DMA_Addr_Translation:master_write -> mm_interconnect_0:Video_In_DMA_Addr_Translation_master_write
	wire  [31:0] video_in_dma_addr_translation_master_writedata;                                        // Video_In_DMA_Addr_Translation:master_writedata -> mm_interconnect_0:Video_In_DMA_Addr_Translation_master_writedata
	wire   [1:0] arm_a9_hps_h2f_axi_master_awburst;                                                     // ARM_A9_HPS:h2f_AWBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awburst
	wire   [3:0] arm_a9_hps_h2f_axi_master_arlen;                                                       // ARM_A9_HPS:h2f_ARLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arlen
	wire   [7:0] arm_a9_hps_h2f_axi_master_wstrb;                                                       // ARM_A9_HPS:h2f_WSTRB -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wstrb
	wire         arm_a9_hps_h2f_axi_master_wready;                                                      // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wready -> ARM_A9_HPS:h2f_WREADY
	wire  [11:0] arm_a9_hps_h2f_axi_master_rid;                                                         // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rid -> ARM_A9_HPS:h2f_RID
	wire         arm_a9_hps_h2f_axi_master_rready;                                                      // ARM_A9_HPS:h2f_RREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rready
	wire   [3:0] arm_a9_hps_h2f_axi_master_awlen;                                                       // ARM_A9_HPS:h2f_AWLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awlen
	wire  [11:0] arm_a9_hps_h2f_axi_master_wid;                                                         // ARM_A9_HPS:h2f_WID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wid
	wire   [3:0] arm_a9_hps_h2f_axi_master_arcache;                                                     // ARM_A9_HPS:h2f_ARCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arcache
	wire         arm_a9_hps_h2f_axi_master_wvalid;                                                      // ARM_A9_HPS:h2f_WVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wvalid
	wire  [29:0] arm_a9_hps_h2f_axi_master_araddr;                                                      // ARM_A9_HPS:h2f_ARADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_araddr
	wire   [2:0] arm_a9_hps_h2f_axi_master_arprot;                                                      // ARM_A9_HPS:h2f_ARPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arprot
	wire   [2:0] arm_a9_hps_h2f_axi_master_awprot;                                                      // ARM_A9_HPS:h2f_AWPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awprot
	wire  [63:0] arm_a9_hps_h2f_axi_master_wdata;                                                       // ARM_A9_HPS:h2f_WDATA -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wdata
	wire         arm_a9_hps_h2f_axi_master_arvalid;                                                     // ARM_A9_HPS:h2f_ARVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arvalid
	wire   [3:0] arm_a9_hps_h2f_axi_master_awcache;                                                     // ARM_A9_HPS:h2f_AWCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awcache
	wire  [11:0] arm_a9_hps_h2f_axi_master_arid;                                                        // ARM_A9_HPS:h2f_ARID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arid
	wire   [1:0] arm_a9_hps_h2f_axi_master_arlock;                                                      // ARM_A9_HPS:h2f_ARLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arlock
	wire   [1:0] arm_a9_hps_h2f_axi_master_awlock;                                                      // ARM_A9_HPS:h2f_AWLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awlock
	wire  [29:0] arm_a9_hps_h2f_axi_master_awaddr;                                                      // ARM_A9_HPS:h2f_AWADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awaddr
	wire   [1:0] arm_a9_hps_h2f_axi_master_bresp;                                                       // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bresp -> ARM_A9_HPS:h2f_BRESP
	wire         arm_a9_hps_h2f_axi_master_arready;                                                     // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arready -> ARM_A9_HPS:h2f_ARREADY
	wire  [63:0] arm_a9_hps_h2f_axi_master_rdata;                                                       // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rdata -> ARM_A9_HPS:h2f_RDATA
	wire         arm_a9_hps_h2f_axi_master_awready;                                                     // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awready -> ARM_A9_HPS:h2f_AWREADY
	wire   [1:0] arm_a9_hps_h2f_axi_master_arburst;                                                     // ARM_A9_HPS:h2f_ARBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arburst
	wire   [2:0] arm_a9_hps_h2f_axi_master_arsize;                                                      // ARM_A9_HPS:h2f_ARSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arsize
	wire         arm_a9_hps_h2f_axi_master_bready;                                                      // ARM_A9_HPS:h2f_BREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bready
	wire         arm_a9_hps_h2f_axi_master_rlast;                                                       // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rlast -> ARM_A9_HPS:h2f_RLAST
	wire         arm_a9_hps_h2f_axi_master_wlast;                                                       // ARM_A9_HPS:h2f_WLAST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wlast
	wire   [1:0] arm_a9_hps_h2f_axi_master_rresp;                                                       // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rresp -> ARM_A9_HPS:h2f_RRESP
	wire  [11:0] arm_a9_hps_h2f_axi_master_awid;                                                        // ARM_A9_HPS:h2f_AWID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awid
	wire  [11:0] arm_a9_hps_h2f_axi_master_bid;                                                         // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bid -> ARM_A9_HPS:h2f_BID
	wire         arm_a9_hps_h2f_axi_master_bvalid;                                                      // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bvalid -> ARM_A9_HPS:h2f_BVALID
	wire   [2:0] arm_a9_hps_h2f_axi_master_awsize;                                                      // ARM_A9_HPS:h2f_AWSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awsize
	wire         arm_a9_hps_h2f_axi_master_awvalid;                                                     // ARM_A9_HPS:h2f_AWVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awvalid
	wire         arm_a9_hps_h2f_axi_master_rvalid;                                                      // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rvalid -> ARM_A9_HPS:h2f_RVALID
	wire         video_in_subsystem_video_in_dma_master_waitrequest;                                    // mm_interconnect_0:Video_In_Subsystem_video_in_dma_master_waitrequest -> Video_In_Subsystem:video_in_dma_master_waitrequest
	wire  [31:0] video_in_subsystem_video_in_dma_master_address;                                        // Video_In_Subsystem:video_in_dma_master_address -> mm_interconnect_0:Video_In_Subsystem_video_in_dma_master_address
	wire         video_in_subsystem_video_in_dma_master_write;                                          // Video_In_Subsystem:video_in_dma_master_write -> mm_interconnect_0:Video_In_Subsystem_video_in_dma_master_write
	wire  [15:0] video_in_subsystem_video_in_dma_master_writedata;                                      // Video_In_Subsystem:video_in_dma_master_writedata -> mm_interconnect_0:Video_In_Subsystem_video_in_dma_master_writedata
	wire  [31:0] nios2_2nd_core_instruction_master_readdata;                                            // mm_interconnect_0:Nios2_2nd_Core_instruction_master_readdata -> Nios2_2nd_Core:i_readdata
	wire         nios2_2nd_core_instruction_master_waitrequest;                                         // mm_interconnect_0:Nios2_2nd_Core_instruction_master_waitrequest -> Nios2_2nd_Core:i_waitrequest
	wire  [27:0] nios2_2nd_core_instruction_master_address;                                             // Nios2_2nd_Core:i_address -> mm_interconnect_0:Nios2_2nd_Core_instruction_master_address
	wire         nios2_2nd_core_instruction_master_read;                                                // Nios2_2nd_Core:i_read -> mm_interconnect_0:Nios2_2nd_Core_instruction_master_read
	wire         nios2_2nd_core_instruction_master_readdatavalid;                                       // mm_interconnect_0:Nios2_2nd_Core_instruction_master_readdatavalid -> Nios2_2nd_Core:i_readdatavalid
	wire  [31:0] nios2_instruction_master_readdata;                                                     // mm_interconnect_0:Nios2_instruction_master_readdata -> Nios2:i_readdata
	wire         nios2_instruction_master_waitrequest;                                                  // mm_interconnect_0:Nios2_instruction_master_waitrequest -> Nios2:i_waitrequest
	wire  [27:0] nios2_instruction_master_address;                                                      // Nios2:i_address -> mm_interconnect_0:Nios2_instruction_master_address
	wire         nios2_instruction_master_read;                                                         // Nios2:i_read -> mm_interconnect_0:Nios2_instruction_master_read
	wire         nios2_instruction_master_readdatavalid;                                                // mm_interconnect_0:Nios2_instruction_master_readdatavalid -> Nios2:i_readdatavalid
	wire         vga_subsystem_pixel_dma_master_waitrequest;                                            // mm_interconnect_0:VGA_Subsystem_pixel_dma_master_waitrequest -> VGA_Subsystem:pixel_dma_master_waitrequest
	wire  [15:0] vga_subsystem_pixel_dma_master_readdata;                                               // mm_interconnect_0:VGA_Subsystem_pixel_dma_master_readdata -> VGA_Subsystem:pixel_dma_master_readdata
	wire  [31:0] vga_subsystem_pixel_dma_master_address;                                                // VGA_Subsystem:pixel_dma_master_address -> mm_interconnect_0:VGA_Subsystem_pixel_dma_master_address
	wire         vga_subsystem_pixel_dma_master_read;                                                   // VGA_Subsystem:pixel_dma_master_read -> mm_interconnect_0:VGA_Subsystem_pixel_dma_master_read
	wire         vga_subsystem_pixel_dma_master_readdatavalid;                                          // mm_interconnect_0:VGA_Subsystem_pixel_dma_master_readdatavalid -> VGA_Subsystem:pixel_dma_master_readdatavalid
	wire         vga_subsystem_pixel_dma_master_lock;                                                   // VGA_Subsystem:pixel_dma_master_lock -> mm_interconnect_0:VGA_Subsystem_pixel_dma_master_lock
	wire  [31:0] pixel_dma_addr_translation_master_readdata;                                            // mm_interconnect_0:Pixel_DMA_Addr_Translation_master_readdata -> Pixel_DMA_Addr_Translation:master_readdata
	wire         pixel_dma_addr_translation_master_waitrequest;                                         // mm_interconnect_0:Pixel_DMA_Addr_Translation_master_waitrequest -> Pixel_DMA_Addr_Translation:master_waitrequest
	wire   [1:0] pixel_dma_addr_translation_master_address;                                             // Pixel_DMA_Addr_Translation:master_address -> mm_interconnect_0:Pixel_DMA_Addr_Translation_master_address
	wire   [3:0] pixel_dma_addr_translation_master_byteenable;                                          // Pixel_DMA_Addr_Translation:master_byteenable -> mm_interconnect_0:Pixel_DMA_Addr_Translation_master_byteenable
	wire         pixel_dma_addr_translation_master_read;                                                // Pixel_DMA_Addr_Translation:master_read -> mm_interconnect_0:Pixel_DMA_Addr_Translation_master_read
	wire         pixel_dma_addr_translation_master_write;                                               // Pixel_DMA_Addr_Translation:master_write -> mm_interconnect_0:Pixel_DMA_Addr_Translation_master_write
	wire  [31:0] pixel_dma_addr_translation_master_writedata;                                           // Pixel_DMA_Addr_Translation:master_writedata -> mm_interconnect_0:Pixel_DMA_Addr_Translation_master_writedata
	wire  [31:0] char_dma_addr_translation_master_readdata;                                             // mm_interconnect_0:Char_DMA_Addr_Translation_master_readdata -> Char_DMA_Addr_Translation:master_readdata
	wire         char_dma_addr_translation_master_waitrequest;                                          // mm_interconnect_0:Char_DMA_Addr_Translation_master_waitrequest -> Char_DMA_Addr_Translation:master_waitrequest
	wire   [1:0] char_dma_addr_translation_master_address;                                              // Char_DMA_Addr_Translation:master_address -> mm_interconnect_0:Char_DMA_Addr_Translation_master_address
	wire   [3:0] char_dma_addr_translation_master_byteenable;                                           // Char_DMA_Addr_Translation:master_byteenable -> mm_interconnect_0:Char_DMA_Addr_Translation_master_byteenable
	wire         char_dma_addr_translation_master_read;                                                 // Char_DMA_Addr_Translation:master_read -> mm_interconnect_0:Char_DMA_Addr_Translation_master_read
	wire         char_dma_addr_translation_master_write;                                                // Char_DMA_Addr_Translation:master_write -> mm_interconnect_0:Char_DMA_Addr_Translation_master_write
	wire  [31:0] char_dma_addr_translation_master_writedata;                                            // Char_DMA_Addr_Translation:master_writedata -> mm_interconnect_0:Char_DMA_Addr_Translation_master_writedata
	wire  [31:0] mm_interconnect_0_adc_adc_slave_readdata;                                              // ADC:readdata -> mm_interconnect_0:ADC_adc_slave_readdata
	wire         mm_interconnect_0_adc_adc_slave_waitrequest;                                           // ADC:waitrequest -> mm_interconnect_0:ADC_adc_slave_waitrequest
	wire   [2:0] mm_interconnect_0_adc_adc_slave_address;                                               // mm_interconnect_0:ADC_adc_slave_address -> ADC:address
	wire         mm_interconnect_0_adc_adc_slave_read;                                                  // mm_interconnect_0:ADC_adc_slave_read -> ADC:read
	wire         mm_interconnect_0_adc_adc_slave_write;                                                 // mm_interconnect_0:ADC_adc_slave_write -> ADC:write
	wire  [31:0] mm_interconnect_0_adc_adc_slave_writedata;                                             // mm_interconnect_0:ADC_adc_slave_writedata -> ADC:writedata
	wire         mm_interconnect_0_audio_subsystem_audio_slave_chipselect;                              // mm_interconnect_0:Audio_Subsystem_audio_slave_chipselect -> Audio_Subsystem:audio_slave_chipselect
	wire  [31:0] mm_interconnect_0_audio_subsystem_audio_slave_readdata;                                // Audio_Subsystem:audio_slave_readdata -> mm_interconnect_0:Audio_Subsystem_audio_slave_readdata
	wire   [1:0] mm_interconnect_0_audio_subsystem_audio_slave_address;                                 // mm_interconnect_0:Audio_Subsystem_audio_slave_address -> Audio_Subsystem:audio_slave_address
	wire         mm_interconnect_0_audio_subsystem_audio_slave_read;                                    // mm_interconnect_0:Audio_Subsystem_audio_slave_read -> Audio_Subsystem:audio_slave_read
	wire         mm_interconnect_0_audio_subsystem_audio_slave_write;                                   // mm_interconnect_0:Audio_Subsystem_audio_slave_write -> Audio_Subsystem:audio_slave_write
	wire  [31:0] mm_interconnect_0_audio_subsystem_audio_slave_writedata;                               // mm_interconnect_0:Audio_Subsystem_audio_slave_writedata -> Audio_Subsystem:audio_slave_writedata
	wire  [31:0] mm_interconnect_0_av_config_avalon_av_config_slave_readdata;                           // AV_Config:readdata -> mm_interconnect_0:AV_Config_avalon_av_config_slave_readdata
	wire         mm_interconnect_0_av_config_avalon_av_config_slave_waitrequest;                        // AV_Config:waitrequest -> mm_interconnect_0:AV_Config_avalon_av_config_slave_waitrequest
	wire   [1:0] mm_interconnect_0_av_config_avalon_av_config_slave_address;                            // mm_interconnect_0:AV_Config_avalon_av_config_slave_address -> AV_Config:address
	wire         mm_interconnect_0_av_config_avalon_av_config_slave_read;                               // mm_interconnect_0:AV_Config_avalon_av_config_slave_read -> AV_Config:read
	wire   [3:0] mm_interconnect_0_av_config_avalon_av_config_slave_byteenable;                         // mm_interconnect_0:AV_Config_avalon_av_config_slave_byteenable -> AV_Config:byteenable
	wire         mm_interconnect_0_av_config_avalon_av_config_slave_write;                              // mm_interconnect_0:AV_Config_avalon_av_config_slave_write -> AV_Config:write
	wire  [31:0] mm_interconnect_0_av_config_avalon_av_config_slave_writedata;                          // mm_interconnect_0:AV_Config_avalon_av_config_slave_writedata -> AV_Config:writedata
	wire         mm_interconnect_0_irda_avalon_irda_slave_chipselect;                                   // mm_interconnect_0:IrDA_avalon_irda_slave_chipselect -> IrDA:chipselect
	wire  [31:0] mm_interconnect_0_irda_avalon_irda_slave_readdata;                                     // IrDA:readdata -> mm_interconnect_0:IrDA_avalon_irda_slave_readdata
	wire   [0:0] mm_interconnect_0_irda_avalon_irda_slave_address;                                      // mm_interconnect_0:IrDA_avalon_irda_slave_address -> IrDA:address
	wire         mm_interconnect_0_irda_avalon_irda_slave_read;                                         // mm_interconnect_0:IrDA_avalon_irda_slave_read -> IrDA:read
	wire   [3:0] mm_interconnect_0_irda_avalon_irda_slave_byteenable;                                   // mm_interconnect_0:IrDA_avalon_irda_slave_byteenable -> IrDA:byteenable
	wire         mm_interconnect_0_irda_avalon_irda_slave_write;                                        // mm_interconnect_0:IrDA_avalon_irda_slave_write -> IrDA:write
	wire  [31:0] mm_interconnect_0_irda_avalon_irda_slave_writedata;                                    // mm_interconnect_0:IrDA_avalon_irda_slave_writedata -> IrDA:writedata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                              // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                                // JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                             // JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                                 // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                                    // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> JTAG_UART:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                                   // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> JTAG_UART:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                               // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	wire         mm_interconnect_0_ps2_port_avalon_ps2_slave_chipselect;                                // mm_interconnect_0:PS2_Port_avalon_ps2_slave_chipselect -> PS2_Port:chipselect
	wire  [31:0] mm_interconnect_0_ps2_port_avalon_ps2_slave_readdata;                                  // PS2_Port:readdata -> mm_interconnect_0:PS2_Port_avalon_ps2_slave_readdata
	wire         mm_interconnect_0_ps2_port_avalon_ps2_slave_waitrequest;                               // PS2_Port:waitrequest -> mm_interconnect_0:PS2_Port_avalon_ps2_slave_waitrequest
	wire   [0:0] mm_interconnect_0_ps2_port_avalon_ps2_slave_address;                                   // mm_interconnect_0:PS2_Port_avalon_ps2_slave_address -> PS2_Port:address
	wire         mm_interconnect_0_ps2_port_avalon_ps2_slave_read;                                      // mm_interconnect_0:PS2_Port_avalon_ps2_slave_read -> PS2_Port:read
	wire   [3:0] mm_interconnect_0_ps2_port_avalon_ps2_slave_byteenable;                                // mm_interconnect_0:PS2_Port_avalon_ps2_slave_byteenable -> PS2_Port:byteenable
	wire         mm_interconnect_0_ps2_port_avalon_ps2_slave_write;                                     // mm_interconnect_0:PS2_Port_avalon_ps2_slave_write -> PS2_Port:write
	wire  [31:0] mm_interconnect_0_ps2_port_avalon_ps2_slave_writedata;                                 // mm_interconnect_0:PS2_Port_avalon_ps2_slave_writedata -> PS2_Port:writedata
	wire         mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_chipselect;                           // mm_interconnect_0:PS2_Port_Dual_avalon_ps2_slave_chipselect -> PS2_Port_Dual:chipselect
	wire  [31:0] mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_readdata;                             // PS2_Port_Dual:readdata -> mm_interconnect_0:PS2_Port_Dual_avalon_ps2_slave_readdata
	wire         mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_waitrequest;                          // PS2_Port_Dual:waitrequest -> mm_interconnect_0:PS2_Port_Dual_avalon_ps2_slave_waitrequest
	wire   [0:0] mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_address;                              // mm_interconnect_0:PS2_Port_Dual_avalon_ps2_slave_address -> PS2_Port_Dual:address
	wire         mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_read;                                 // mm_interconnect_0:PS2_Port_Dual_avalon_ps2_slave_read -> PS2_Port_Dual:read
	wire   [3:0] mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_byteenable;                           // mm_interconnect_0:PS2_Port_Dual_avalon_ps2_slave_byteenable -> PS2_Port_Dual:byteenable
	wire         mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_write;                                // mm_interconnect_0:PS2_Port_Dual_avalon_ps2_slave_write -> PS2_Port_Dual:write
	wire  [31:0] mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_writedata;                            // mm_interconnect_0:PS2_Port_Dual_avalon_ps2_slave_writedata -> PS2_Port_Dual:writedata
	wire  [31:0] mm_interconnect_0_vga_subsystem_char_buffer_control_slave_readdata;                    // VGA_Subsystem:char_buffer_control_slave_readdata -> mm_interconnect_0:VGA_Subsystem_char_buffer_control_slave_readdata
	wire   [1:0] mm_interconnect_0_vga_subsystem_char_buffer_control_slave_address;                     // mm_interconnect_0:VGA_Subsystem_char_buffer_control_slave_address -> VGA_Subsystem:char_buffer_control_slave_address
	wire         mm_interconnect_0_vga_subsystem_char_buffer_control_slave_read;                        // mm_interconnect_0:VGA_Subsystem_char_buffer_control_slave_read -> VGA_Subsystem:char_buffer_control_slave_read
	wire   [3:0] mm_interconnect_0_vga_subsystem_char_buffer_control_slave_byteenable;                  // mm_interconnect_0:VGA_Subsystem_char_buffer_control_slave_byteenable -> VGA_Subsystem:char_buffer_control_slave_byteenable
	wire         mm_interconnect_0_vga_subsystem_char_buffer_control_slave_write;                       // mm_interconnect_0:VGA_Subsystem_char_buffer_control_slave_write -> VGA_Subsystem:char_buffer_control_slave_write
	wire  [31:0] mm_interconnect_0_vga_subsystem_char_buffer_control_slave_writedata;                   // mm_interconnect_0:VGA_Subsystem_char_buffer_control_slave_writedata -> VGA_Subsystem:char_buffer_control_slave_writedata
	wire         mm_interconnect_0_vga_subsystem_char_buffer_slave_chipselect;                          // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_chipselect -> VGA_Subsystem:char_buffer_slave_chipselect
	wire  [31:0] mm_interconnect_0_vga_subsystem_char_buffer_slave_readdata;                            // VGA_Subsystem:char_buffer_slave_readdata -> mm_interconnect_0:VGA_Subsystem_char_buffer_slave_readdata
	wire  [10:0] mm_interconnect_0_vga_subsystem_char_buffer_slave_address;                             // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_address -> VGA_Subsystem:char_buffer_slave_address
	wire   [3:0] mm_interconnect_0_vga_subsystem_char_buffer_slave_byteenable;                          // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_byteenable -> VGA_Subsystem:char_buffer_slave_byteenable
	wire         mm_interconnect_0_vga_subsystem_char_buffer_slave_write;                               // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_write -> VGA_Subsystem:char_buffer_slave_write
	wire  [31:0] mm_interconnect_0_vga_subsystem_char_buffer_slave_writedata;                           // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_writedata -> VGA_Subsystem:char_buffer_slave_writedata
	wire         mm_interconnect_0_vga_subsystem_char_buffer_slave_clken;                               // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_clken -> VGA_Subsystem:char_buffer_slave_clken
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                                        // SysID:readdata -> mm_interconnect_0:SysID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                                         // mm_interconnect_0:SysID_control_slave_address -> SysID:address
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;                                      // Nios2:debug_mem_slave_readdata -> mm_interconnect_0:Nios2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;                                   // Nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:Nios2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;                                   // mm_interconnect_0:Nios2_debug_mem_slave_debugaccess -> Nios2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;                                       // mm_interconnect_0:Nios2_debug_mem_slave_address -> Nios2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;                                          // mm_interconnect_0:Nios2_debug_mem_slave_read -> Nios2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;                                    // mm_interconnect_0:Nios2_debug_mem_slave_byteenable -> Nios2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;                                         // mm_interconnect_0:Nios2_debug_mem_slave_write -> Nios2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;                                     // mm_interconnect_0:Nios2_debug_mem_slave_writedata -> Nios2:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_readdata;                      // VGA_Subsystem:pixel_dma_control_slave_readdata -> mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_readdata
	wire   [1:0] mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_address;                       // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_address -> VGA_Subsystem:pixel_dma_control_slave_address
	wire         mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_read;                          // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_read -> VGA_Subsystem:pixel_dma_control_slave_read
	wire   [3:0] mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_byteenable;                    // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_byteenable -> VGA_Subsystem:pixel_dma_control_slave_byteenable
	wire         mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_write;                         // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_write -> VGA_Subsystem:pixel_dma_control_slave_write
	wire  [31:0] mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_writedata;                     // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_writedata -> VGA_Subsystem:pixel_dma_control_slave_writedata
	wire  [31:0] mm_interconnect_0_vga_subsystem_rgb_slave_readdata;                                    // VGA_Subsystem:rgb_slave_readdata -> mm_interconnect_0:VGA_Subsystem_rgb_slave_readdata
	wire         mm_interconnect_0_vga_subsystem_rgb_slave_read;                                        // mm_interconnect_0:VGA_Subsystem_rgb_slave_read -> VGA_Subsystem:rgb_slave_read
	wire         mm_interconnect_0_sdram_s1_chipselect;                                                 // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                                   // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                                // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                                    // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                                       // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                                 // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                              // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                                      // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                                  // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire         mm_interconnect_0_onchip_sram_s1_chipselect;                                           // mm_interconnect_0:Onchip_SRAM_s1_chipselect -> Onchip_SRAM:chipselect
	wire  [31:0] mm_interconnect_0_onchip_sram_s1_readdata;                                             // Onchip_SRAM:readdata -> mm_interconnect_0:Onchip_SRAM_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_sram_s1_address;                                              // mm_interconnect_0:Onchip_SRAM_s1_address -> Onchip_SRAM:address
	wire   [3:0] mm_interconnect_0_onchip_sram_s1_byteenable;                                           // mm_interconnect_0:Onchip_SRAM_s1_byteenable -> Onchip_SRAM:byteenable
	wire         mm_interconnect_0_onchip_sram_s1_write;                                                // mm_interconnect_0:Onchip_SRAM_s1_write -> Onchip_SRAM:write
	wire  [31:0] mm_interconnect_0_onchip_sram_s1_writedata;                                            // mm_interconnect_0:Onchip_SRAM_s1_writedata -> Onchip_SRAM:writedata
	wire         mm_interconnect_0_onchip_sram_s1_clken;                                                // mm_interconnect_0:Onchip_SRAM_s1_clken -> Onchip_SRAM:clken
	wire         mm_interconnect_0_leds_s1_chipselect;                                                  // mm_interconnect_0:LEDs_s1_chipselect -> LEDs:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                                                    // LEDs:readdata -> mm_interconnect_0:LEDs_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                                                     // mm_interconnect_0:LEDs_s1_address -> LEDs:address
	wire         mm_interconnect_0_leds_s1_write;                                                       // mm_interconnect_0:LEDs_s1_write -> LEDs:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                                                   // mm_interconnect_0:LEDs_s1_writedata -> LEDs:writedata
	wire         mm_interconnect_0_hex3_hex0_s1_chipselect;                                             // mm_interconnect_0:HEX3_HEX0_s1_chipselect -> HEX3_HEX0:chipselect
	wire  [31:0] mm_interconnect_0_hex3_hex0_s1_readdata;                                               // HEX3_HEX0:readdata -> mm_interconnect_0:HEX3_HEX0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex3_hex0_s1_address;                                                // mm_interconnect_0:HEX3_HEX0_s1_address -> HEX3_HEX0:address
	wire         mm_interconnect_0_hex3_hex0_s1_write;                                                  // mm_interconnect_0:HEX3_HEX0_s1_write -> HEX3_HEX0:write_n
	wire  [31:0] mm_interconnect_0_hex3_hex0_s1_writedata;                                              // mm_interconnect_0:HEX3_HEX0_s1_writedata -> HEX3_HEX0:writedata
	wire         mm_interconnect_0_hex5_hex4_s1_chipselect;                                             // mm_interconnect_0:HEX5_HEX4_s1_chipselect -> HEX5_HEX4:chipselect
	wire  [31:0] mm_interconnect_0_hex5_hex4_s1_readdata;                                               // HEX5_HEX4:readdata -> mm_interconnect_0:HEX5_HEX4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex5_hex4_s1_address;                                                // mm_interconnect_0:HEX5_HEX4_s1_address -> HEX5_HEX4:address
	wire         mm_interconnect_0_hex5_hex4_s1_write;                                                  // mm_interconnect_0:HEX5_HEX4_s1_write -> HEX5_HEX4:write_n
	wire  [31:0] mm_interconnect_0_hex5_hex4_s1_writedata;                                              // mm_interconnect_0:HEX5_HEX4_s1_writedata -> HEX5_HEX4:writedata
	wire  [31:0] mm_interconnect_0_slider_switches_s1_readdata;                                         // Slider_Switches:readdata -> mm_interconnect_0:Slider_Switches_s1_readdata
	wire   [1:0] mm_interconnect_0_slider_switches_s1_address;                                          // mm_interconnect_0:Slider_Switches_s1_address -> Slider_Switches:address
	wire         mm_interconnect_0_pushbuttons_s1_chipselect;                                           // mm_interconnect_0:Pushbuttons_s1_chipselect -> Pushbuttons:chipselect
	wire  [31:0] mm_interconnect_0_pushbuttons_s1_readdata;                                             // Pushbuttons:readdata -> mm_interconnect_0:Pushbuttons_s1_readdata
	wire   [1:0] mm_interconnect_0_pushbuttons_s1_address;                                              // mm_interconnect_0:Pushbuttons_s1_address -> Pushbuttons:address
	wire         mm_interconnect_0_pushbuttons_s1_write;                                                // mm_interconnect_0:Pushbuttons_s1_write -> Pushbuttons:write_n
	wire  [31:0] mm_interconnect_0_pushbuttons_s1_writedata;                                            // mm_interconnect_0:Pushbuttons_s1_writedata -> Pushbuttons:writedata
	wire         mm_interconnect_0_expansion_jp1_s1_chipselect;                                         // mm_interconnect_0:Expansion_JP1_s1_chipselect -> Expansion_JP1:chipselect
	wire  [31:0] mm_interconnect_0_expansion_jp1_s1_readdata;                                           // Expansion_JP1:readdata -> mm_interconnect_0:Expansion_JP1_s1_readdata
	wire   [1:0] mm_interconnect_0_expansion_jp1_s1_address;                                            // mm_interconnect_0:Expansion_JP1_s1_address -> Expansion_JP1:address
	wire         mm_interconnect_0_expansion_jp1_s1_write;                                              // mm_interconnect_0:Expansion_JP1_s1_write -> Expansion_JP1:write_n
	wire  [31:0] mm_interconnect_0_expansion_jp1_s1_writedata;                                          // mm_interconnect_0:Expansion_JP1_s1_writedata -> Expansion_JP1:writedata
	wire         mm_interconnect_0_interval_timer_s1_chipselect;                                        // mm_interconnect_0:Interval_Timer_s1_chipselect -> Interval_Timer:chipselect
	wire  [15:0] mm_interconnect_0_interval_timer_s1_readdata;                                          // Interval_Timer:readdata -> mm_interconnect_0:Interval_Timer_s1_readdata
	wire   [2:0] mm_interconnect_0_interval_timer_s1_address;                                           // mm_interconnect_0:Interval_Timer_s1_address -> Interval_Timer:address
	wire         mm_interconnect_0_interval_timer_s1_write;                                             // mm_interconnect_0:Interval_Timer_s1_write -> Interval_Timer:write_n
	wire  [15:0] mm_interconnect_0_interval_timer_s1_writedata;                                         // mm_interconnect_0:Interval_Timer_s1_writedata -> Interval_Timer:writedata
	wire         mm_interconnect_0_interval_timer_2_s1_chipselect;                                      // mm_interconnect_0:Interval_Timer_2_s1_chipselect -> Interval_Timer_2:chipselect
	wire  [15:0] mm_interconnect_0_interval_timer_2_s1_readdata;                                        // Interval_Timer_2:readdata -> mm_interconnect_0:Interval_Timer_2_s1_readdata
	wire   [2:0] mm_interconnect_0_interval_timer_2_s1_address;                                         // mm_interconnect_0:Interval_Timer_2_s1_address -> Interval_Timer_2:address
	wire         mm_interconnect_0_interval_timer_2_s1_write;                                           // mm_interconnect_0:Interval_Timer_2_s1_write -> Interval_Timer_2:write_n
	wire  [15:0] mm_interconnect_0_interval_timer_2_s1_writedata;                                       // mm_interconnect_0:Interval_Timer_2_s1_writedata -> Interval_Timer_2:writedata
	wire  [31:0] mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_readdata;              // Video_In_Subsystem:video_in_dma_control_slave_readdata -> mm_interconnect_0:Video_In_Subsystem_video_in_dma_control_slave_readdata
	wire   [1:0] mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_address;               // mm_interconnect_0:Video_In_Subsystem_video_in_dma_control_slave_address -> Video_In_Subsystem:video_in_dma_control_slave_address
	wire         mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_read;                  // mm_interconnect_0:Video_In_Subsystem_video_in_dma_control_slave_read -> Video_In_Subsystem:video_in_dma_control_slave_read
	wire   [3:0] mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_byteenable;            // mm_interconnect_0:Video_In_Subsystem_video_in_dma_control_slave_byteenable -> Video_In_Subsystem:video_in_dma_control_slave_byteenable
	wire         mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_write;                 // mm_interconnect_0:Video_In_Subsystem_video_in_dma_control_slave_write -> Video_In_Subsystem:video_in_dma_control_slave_write
	wire  [31:0] mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_writedata;             // mm_interconnect_0:Video_In_Subsystem_video_in_dma_control_slave_writedata -> Video_In_Subsystem:video_in_dma_control_slave_writedata
	wire         mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_chipselect; // mm_interconnect_0:Video_In_Subsystem_video_in_edge_detection_control_slave_chipselect -> Video_In_Subsystem:video_in_edge_detection_control_slave_chipselect
	wire  [31:0] mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_readdata;   // Video_In_Subsystem:video_in_edge_detection_control_slave_readdata -> mm_interconnect_0:Video_In_Subsystem_video_in_edge_detection_control_slave_readdata
	wire   [1:0] mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_address;    // mm_interconnect_0:Video_In_Subsystem_video_in_edge_detection_control_slave_address -> Video_In_Subsystem:video_in_edge_detection_control_slave_address
	wire         mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_write;      // mm_interconnect_0:Video_In_Subsystem_video_in_edge_detection_control_slave_write -> Video_In_Subsystem:video_in_edge_detection_control_slave_write_n
	wire  [31:0] mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_writedata;  // mm_interconnect_0:Video_In_Subsystem_video_in_edge_detection_control_slave_writedata -> Video_In_Subsystem:video_in_edge_detection_control_slave_writedata
	wire  [31:0] mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_readdata;                     // F2H_Mem_Window_00000000:avs_s0_readdata -> mm_interconnect_0:F2H_Mem_Window_00000000_windowed_slave_readdata
	wire         mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_waitrequest;                  // F2H_Mem_Window_00000000:avs_s0_waitrequest -> mm_interconnect_0:F2H_Mem_Window_00000000_windowed_slave_waitrequest
	wire  [27:0] mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_address;                      // mm_interconnect_0:F2H_Mem_Window_00000000_windowed_slave_address -> F2H_Mem_Window_00000000:avs_s0_address
	wire         mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_read;                         // mm_interconnect_0:F2H_Mem_Window_00000000_windowed_slave_read -> F2H_Mem_Window_00000000:avs_s0_read
	wire   [3:0] mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_byteenable;                   // mm_interconnect_0:F2H_Mem_Window_00000000_windowed_slave_byteenable -> F2H_Mem_Window_00000000:avs_s0_byteenable
	wire         mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_readdatavalid;                // F2H_Mem_Window_00000000:avs_s0_readdatavalid -> mm_interconnect_0:F2H_Mem_Window_00000000_windowed_slave_readdatavalid
	wire         mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_write;                        // mm_interconnect_0:F2H_Mem_Window_00000000_windowed_slave_write -> F2H_Mem_Window_00000000:avs_s0_write
	wire  [31:0] mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_writedata;                    // mm_interconnect_0:F2H_Mem_Window_00000000_windowed_slave_writedata -> F2H_Mem_Window_00000000:avs_s0_writedata
	wire   [0:0] mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_burstcount;                   // mm_interconnect_0:F2H_Mem_Window_00000000_windowed_slave_burstcount -> F2H_Mem_Window_00000000:avs_s0_burstcount
	wire  [31:0] mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_readdata;                     // F2H_Mem_Window_FF600000:avs_s0_readdata -> mm_interconnect_0:F2H_Mem_Window_FF600000_windowed_slave_readdata
	wire         mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_waitrequest;                  // F2H_Mem_Window_FF600000:avs_s0_waitrequest -> mm_interconnect_0:F2H_Mem_Window_FF600000_windowed_slave_waitrequest
	wire  [18:0] mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_address;                      // mm_interconnect_0:F2H_Mem_Window_FF600000_windowed_slave_address -> F2H_Mem_Window_FF600000:avs_s0_address
	wire         mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_read;                         // mm_interconnect_0:F2H_Mem_Window_FF600000_windowed_slave_read -> F2H_Mem_Window_FF600000:avs_s0_read
	wire   [3:0] mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_byteenable;                   // mm_interconnect_0:F2H_Mem_Window_FF600000_windowed_slave_byteenable -> F2H_Mem_Window_FF600000:avs_s0_byteenable
	wire         mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_readdatavalid;                // F2H_Mem_Window_FF600000:avs_s0_readdatavalid -> mm_interconnect_0:F2H_Mem_Window_FF600000_windowed_slave_readdatavalid
	wire         mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_write;                        // mm_interconnect_0:F2H_Mem_Window_FF600000_windowed_slave_write -> F2H_Mem_Window_FF600000:avs_s0_write
	wire  [31:0] mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_writedata;                    // mm_interconnect_0:F2H_Mem_Window_FF600000_windowed_slave_writedata -> F2H_Mem_Window_FF600000:avs_s0_writedata
	wire   [0:0] mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_burstcount;                   // mm_interconnect_0:F2H_Mem_Window_FF600000_windowed_slave_burstcount -> F2H_Mem_Window_FF600000:avs_s0_burstcount
	wire  [31:0] mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_readdata;                     // F2H_Mem_Window_FF800000:avs_s0_readdata -> mm_interconnect_0:F2H_Mem_Window_FF800000_windowed_slave_readdata
	wire         mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_waitrequest;                  // F2H_Mem_Window_FF800000:avs_s0_waitrequest -> mm_interconnect_0:F2H_Mem_Window_FF800000_windowed_slave_waitrequest
	wire  [20:0] mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_address;                      // mm_interconnect_0:F2H_Mem_Window_FF800000_windowed_slave_address -> F2H_Mem_Window_FF800000:avs_s0_address
	wire         mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_read;                         // mm_interconnect_0:F2H_Mem_Window_FF800000_windowed_slave_read -> F2H_Mem_Window_FF800000:avs_s0_read
	wire   [3:0] mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_byteenable;                   // mm_interconnect_0:F2H_Mem_Window_FF800000_windowed_slave_byteenable -> F2H_Mem_Window_FF800000:avs_s0_byteenable
	wire         mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_readdatavalid;                // F2H_Mem_Window_FF800000:avs_s0_readdatavalid -> mm_interconnect_0:F2H_Mem_Window_FF800000_windowed_slave_readdatavalid
	wire         mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_write;                        // mm_interconnect_0:F2H_Mem_Window_FF800000_windowed_slave_write -> F2H_Mem_Window_FF800000:avs_s0_write
	wire  [31:0] mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_writedata;                    // mm_interconnect_0:F2H_Mem_Window_FF800000_windowed_slave_writedata -> F2H_Mem_Window_FF800000:avs_s0_writedata
	wire   [0:0] mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_burstcount;                   // mm_interconnect_0:F2H_Mem_Window_FF800000_windowed_slave_burstcount -> F2H_Mem_Window_FF800000:avs_s0_burstcount
	wire         mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_chipselect;                     // mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_chipselect -> JTAG_UART_2nd_Core:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_readdata;                       // JTAG_UART_2nd_Core:av_readdata -> mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_waitrequest;                    // JTAG_UART_2nd_Core:av_waitrequest -> mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_address;                        // mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_address -> JTAG_UART_2nd_Core:av_address
	wire         mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read;                           // mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_read -> JTAG_UART_2nd_Core:av_read_n
	wire         mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write;                          // mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_write -> JTAG_UART_2nd_Core:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_writedata;                      // mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_writedata -> JTAG_UART_2nd_Core:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_2nd_core_debug_mem_slave_readdata;                             // Nios2_2nd_Core:debug_mem_slave_readdata -> mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_2nd_core_debug_mem_slave_waitrequest;                          // Nios2_2nd_Core:debug_mem_slave_waitrequest -> mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_2nd_core_debug_mem_slave_debugaccess;                          // mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_debugaccess -> Nios2_2nd_Core:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_2nd_core_debug_mem_slave_address;                              // mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_address -> Nios2_2nd_Core:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_2nd_core_debug_mem_slave_read;                                 // mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_read -> Nios2_2nd_Core:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_2nd_core_debug_mem_slave_byteenable;                           // mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_byteenable -> Nios2_2nd_Core:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_2nd_core_debug_mem_slave_write;                                // mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_write -> Nios2_2nd_Core:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_2nd_core_debug_mem_slave_writedata;                            // mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_writedata -> Nios2_2nd_Core:debug_mem_slave_writedata
	wire         mm_interconnect_0_interval_timer_2nd_core_s1_chipselect;                               // mm_interconnect_0:Interval_Timer_2nd_Core_s1_chipselect -> Interval_Timer_2nd_Core:chipselect
	wire  [15:0] mm_interconnect_0_interval_timer_2nd_core_s1_readdata;                                 // Interval_Timer_2nd_Core:readdata -> mm_interconnect_0:Interval_Timer_2nd_Core_s1_readdata
	wire   [2:0] mm_interconnect_0_interval_timer_2nd_core_s1_address;                                  // mm_interconnect_0:Interval_Timer_2nd_Core_s1_address -> Interval_Timer_2nd_Core:address
	wire         mm_interconnect_0_interval_timer_2nd_core_s1_write;                                    // mm_interconnect_0:Interval_Timer_2nd_Core_s1_write -> Interval_Timer_2nd_Core:write_n
	wire  [15:0] mm_interconnect_0_interval_timer_2nd_core_s1_writedata;                                // mm_interconnect_0:Interval_Timer_2nd_Core_s1_writedata -> Interval_Timer_2nd_Core:writedata
	wire         mm_interconnect_0_interval_timer_2nd_core_2_s1_chipselect;                             // mm_interconnect_0:Interval_Timer_2nd_Core_2_s1_chipselect -> Interval_Timer_2nd_Core_2:chipselect
	wire  [15:0] mm_interconnect_0_interval_timer_2nd_core_2_s1_readdata;                               // Interval_Timer_2nd_Core_2:readdata -> mm_interconnect_0:Interval_Timer_2nd_Core_2_s1_readdata
	wire   [2:0] mm_interconnect_0_interval_timer_2nd_core_2_s1_address;                                // mm_interconnect_0:Interval_Timer_2nd_Core_2_s1_address -> Interval_Timer_2nd_Core_2:address
	wire         mm_interconnect_0_interval_timer_2nd_core_2_s1_write;                                  // mm_interconnect_0:Interval_Timer_2nd_Core_2_s1_write -> Interval_Timer_2nd_Core_2:write_n
	wire  [15:0] mm_interconnect_0_interval_timer_2nd_core_2_s1_writedata;                              // mm_interconnect_0:Interval_Timer_2nd_Core_2_s1_writedata -> Interval_Timer_2nd_Core_2:writedata
	wire         mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_chipselect;                    // mm_interconnect_0:JTAG_UART_for_ARM_0_avalon_jtag_slave_chipselect -> JTAG_UART_for_ARM_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_readdata;                      // JTAG_UART_for_ARM_0:av_readdata -> mm_interconnect_0:JTAG_UART_for_ARM_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_waitrequest;                   // JTAG_UART_for_ARM_0:av_waitrequest -> mm_interconnect_0:JTAG_UART_for_ARM_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_address;                       // mm_interconnect_0:JTAG_UART_for_ARM_0_avalon_jtag_slave_address -> JTAG_UART_for_ARM_0:av_address
	wire         mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_read;                          // mm_interconnect_0:JTAG_UART_for_ARM_0_avalon_jtag_slave_read -> JTAG_UART_for_ARM_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_write;                         // mm_interconnect_0:JTAG_UART_for_ARM_0_avalon_jtag_slave_write -> JTAG_UART_for_ARM_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_writedata;                     // mm_interconnect_0:JTAG_UART_for_ARM_0_avalon_jtag_slave_writedata -> JTAG_UART_for_ARM_0:av_writedata
	wire         mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_chipselect;                    // mm_interconnect_0:JTAG_UART_for_ARM_1_avalon_jtag_slave_chipselect -> JTAG_UART_for_ARM_1:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_readdata;                      // JTAG_UART_for_ARM_1:av_readdata -> mm_interconnect_0:JTAG_UART_for_ARM_1_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_waitrequest;                   // JTAG_UART_for_ARM_1:av_waitrequest -> mm_interconnect_0:JTAG_UART_for_ARM_1_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_address;                       // mm_interconnect_0:JTAG_UART_for_ARM_1_avalon_jtag_slave_address -> JTAG_UART_for_ARM_1:av_address
	wire         mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_read;                          // mm_interconnect_0:JTAG_UART_for_ARM_1_avalon_jtag_slave_read -> JTAG_UART_for_ARM_1:av_read_n
	wire         mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_write;                         // mm_interconnect_0:JTAG_UART_for_ARM_1_avalon_jtag_slave_write -> JTAG_UART_for_ARM_1:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_writedata;                     // mm_interconnect_0:JTAG_UART_for_ARM_1_avalon_jtag_slave_writedata -> JTAG_UART_for_ARM_1:av_writedata
	wire  [31:0] mm_interconnect_0_pixel_dma_addr_translation_slave_readdata;                           // Pixel_DMA_Addr_Translation:slave_readdata -> mm_interconnect_0:Pixel_DMA_Addr_Translation_slave_readdata
	wire         mm_interconnect_0_pixel_dma_addr_translation_slave_waitrequest;                        // Pixel_DMA_Addr_Translation:slave_waitrequest -> mm_interconnect_0:Pixel_DMA_Addr_Translation_slave_waitrequest
	wire   [1:0] mm_interconnect_0_pixel_dma_addr_translation_slave_address;                            // mm_interconnect_0:Pixel_DMA_Addr_Translation_slave_address -> Pixel_DMA_Addr_Translation:slave_address
	wire         mm_interconnect_0_pixel_dma_addr_translation_slave_read;                               // mm_interconnect_0:Pixel_DMA_Addr_Translation_slave_read -> Pixel_DMA_Addr_Translation:slave_read
	wire   [3:0] mm_interconnect_0_pixel_dma_addr_translation_slave_byteenable;                         // mm_interconnect_0:Pixel_DMA_Addr_Translation_slave_byteenable -> Pixel_DMA_Addr_Translation:slave_byteenable
	wire         mm_interconnect_0_pixel_dma_addr_translation_slave_write;                              // mm_interconnect_0:Pixel_DMA_Addr_Translation_slave_write -> Pixel_DMA_Addr_Translation:slave_write
	wire  [31:0] mm_interconnect_0_pixel_dma_addr_translation_slave_writedata;                          // mm_interconnect_0:Pixel_DMA_Addr_Translation_slave_writedata -> Pixel_DMA_Addr_Translation:slave_writedata
	wire  [31:0] mm_interconnect_0_char_dma_addr_translation_slave_readdata;                            // Char_DMA_Addr_Translation:slave_readdata -> mm_interconnect_0:Char_DMA_Addr_Translation_slave_readdata
	wire         mm_interconnect_0_char_dma_addr_translation_slave_waitrequest;                         // Char_DMA_Addr_Translation:slave_waitrequest -> mm_interconnect_0:Char_DMA_Addr_Translation_slave_waitrequest
	wire   [1:0] mm_interconnect_0_char_dma_addr_translation_slave_address;                             // mm_interconnect_0:Char_DMA_Addr_Translation_slave_address -> Char_DMA_Addr_Translation:slave_address
	wire         mm_interconnect_0_char_dma_addr_translation_slave_read;                                // mm_interconnect_0:Char_DMA_Addr_Translation_slave_read -> Char_DMA_Addr_Translation:slave_read
	wire   [3:0] mm_interconnect_0_char_dma_addr_translation_slave_byteenable;                          // mm_interconnect_0:Char_DMA_Addr_Translation_slave_byteenable -> Char_DMA_Addr_Translation:slave_byteenable
	wire         mm_interconnect_0_char_dma_addr_translation_slave_write;                               // mm_interconnect_0:Char_DMA_Addr_Translation_slave_write -> Char_DMA_Addr_Translation:slave_write
	wire  [31:0] mm_interconnect_0_char_dma_addr_translation_slave_writedata;                           // mm_interconnect_0:Char_DMA_Addr_Translation_slave_writedata -> Char_DMA_Addr_Translation:slave_writedata
	wire  [31:0] mm_interconnect_0_video_in_dma_addr_translation_slave_readdata;                        // Video_In_DMA_Addr_Translation:slave_readdata -> mm_interconnect_0:Video_In_DMA_Addr_Translation_slave_readdata
	wire         mm_interconnect_0_video_in_dma_addr_translation_slave_waitrequest;                     // Video_In_DMA_Addr_Translation:slave_waitrequest -> mm_interconnect_0:Video_In_DMA_Addr_Translation_slave_waitrequest
	wire   [1:0] mm_interconnect_0_video_in_dma_addr_translation_slave_address;                         // mm_interconnect_0:Video_In_DMA_Addr_Translation_slave_address -> Video_In_DMA_Addr_Translation:slave_address
	wire         mm_interconnect_0_video_in_dma_addr_translation_slave_read;                            // mm_interconnect_0:Video_In_DMA_Addr_Translation_slave_read -> Video_In_DMA_Addr_Translation:slave_read
	wire   [3:0] mm_interconnect_0_video_in_dma_addr_translation_slave_byteenable;                      // mm_interconnect_0:Video_In_DMA_Addr_Translation_slave_byteenable -> Video_In_DMA_Addr_Translation:slave_byteenable
	wire         mm_interconnect_0_video_in_dma_addr_translation_slave_write;                           // mm_interconnect_0:Video_In_DMA_Addr_Translation_slave_write -> Video_In_DMA_Addr_Translation:slave_write
	wire  [31:0] mm_interconnect_0_video_in_dma_addr_translation_slave_writedata;                       // mm_interconnect_0:Video_In_DMA_Addr_Translation_slave_writedata -> Video_In_DMA_Addr_Translation:slave_writedata
	wire         mm_interconnect_0_onchip_sram_s2_chipselect;                                           // mm_interconnect_0:Onchip_SRAM_s2_chipselect -> Onchip_SRAM:chipselect2
	wire  [31:0] mm_interconnect_0_onchip_sram_s2_readdata;                                             // Onchip_SRAM:readdata2 -> mm_interconnect_0:Onchip_SRAM_s2_readdata
	wire  [15:0] mm_interconnect_0_onchip_sram_s2_address;                                              // mm_interconnect_0:Onchip_SRAM_s2_address -> Onchip_SRAM:address2
	wire   [3:0] mm_interconnect_0_onchip_sram_s2_byteenable;                                           // mm_interconnect_0:Onchip_SRAM_s2_byteenable -> Onchip_SRAM:byteenable2
	wire         mm_interconnect_0_onchip_sram_s2_write;                                                // mm_interconnect_0:Onchip_SRAM_s2_write -> Onchip_SRAM:write2
	wire  [31:0] mm_interconnect_0_onchip_sram_s2_writedata;                                            // mm_interconnect_0:Onchip_SRAM_s2_writedata -> Onchip_SRAM:writedata2
	wire         mm_interconnect_0_onchip_sram_s2_clken;                                                // mm_interconnect_0:Onchip_SRAM_s2_clken -> Onchip_SRAM:clken2
	wire         f2h_mem_window_00000000_expanded_master_waitrequest;                                   // mm_interconnect_1:F2H_Mem_Window_00000000_expanded_master_waitrequest -> F2H_Mem_Window_00000000:avm_m0_waitrequest
	wire  [31:0] f2h_mem_window_00000000_expanded_master_readdata;                                      // mm_interconnect_1:F2H_Mem_Window_00000000_expanded_master_readdata -> F2H_Mem_Window_00000000:avm_m0_readdata
	wire  [31:0] f2h_mem_window_00000000_expanded_master_address;                                       // F2H_Mem_Window_00000000:avm_m0_address -> mm_interconnect_1:F2H_Mem_Window_00000000_expanded_master_address
	wire         f2h_mem_window_00000000_expanded_master_read;                                          // F2H_Mem_Window_00000000:avm_m0_read -> mm_interconnect_1:F2H_Mem_Window_00000000_expanded_master_read
	wire   [3:0] f2h_mem_window_00000000_expanded_master_byteenable;                                    // F2H_Mem_Window_00000000:avm_m0_byteenable -> mm_interconnect_1:F2H_Mem_Window_00000000_expanded_master_byteenable
	wire         f2h_mem_window_00000000_expanded_master_readdatavalid;                                 // mm_interconnect_1:F2H_Mem_Window_00000000_expanded_master_readdatavalid -> F2H_Mem_Window_00000000:avm_m0_readdatavalid
	wire         f2h_mem_window_00000000_expanded_master_write;                                         // F2H_Mem_Window_00000000:avm_m0_write -> mm_interconnect_1:F2H_Mem_Window_00000000_expanded_master_write
	wire  [31:0] f2h_mem_window_00000000_expanded_master_writedata;                                     // F2H_Mem_Window_00000000:avm_m0_writedata -> mm_interconnect_1:F2H_Mem_Window_00000000_expanded_master_writedata
	wire   [0:0] f2h_mem_window_00000000_expanded_master_burstcount;                                    // F2H_Mem_Window_00000000:avm_m0_burstcount -> mm_interconnect_1:F2H_Mem_Window_00000000_expanded_master_burstcount
	wire         f2h_mem_window_ff600000_expanded_master_waitrequest;                                   // mm_interconnect_1:F2H_Mem_Window_FF600000_expanded_master_waitrequest -> F2H_Mem_Window_FF600000:avm_m0_waitrequest
	wire  [31:0] f2h_mem_window_ff600000_expanded_master_readdata;                                      // mm_interconnect_1:F2H_Mem_Window_FF600000_expanded_master_readdata -> F2H_Mem_Window_FF600000:avm_m0_readdata
	wire  [31:0] f2h_mem_window_ff600000_expanded_master_address;                                       // F2H_Mem_Window_FF600000:avm_m0_address -> mm_interconnect_1:F2H_Mem_Window_FF600000_expanded_master_address
	wire         f2h_mem_window_ff600000_expanded_master_read;                                          // F2H_Mem_Window_FF600000:avm_m0_read -> mm_interconnect_1:F2H_Mem_Window_FF600000_expanded_master_read
	wire   [3:0] f2h_mem_window_ff600000_expanded_master_byteenable;                                    // F2H_Mem_Window_FF600000:avm_m0_byteenable -> mm_interconnect_1:F2H_Mem_Window_FF600000_expanded_master_byteenable
	wire         f2h_mem_window_ff600000_expanded_master_readdatavalid;                                 // mm_interconnect_1:F2H_Mem_Window_FF600000_expanded_master_readdatavalid -> F2H_Mem_Window_FF600000:avm_m0_readdatavalid
	wire         f2h_mem_window_ff600000_expanded_master_write;                                         // F2H_Mem_Window_FF600000:avm_m0_write -> mm_interconnect_1:F2H_Mem_Window_FF600000_expanded_master_write
	wire  [31:0] f2h_mem_window_ff600000_expanded_master_writedata;                                     // F2H_Mem_Window_FF600000:avm_m0_writedata -> mm_interconnect_1:F2H_Mem_Window_FF600000_expanded_master_writedata
	wire   [0:0] f2h_mem_window_ff600000_expanded_master_burstcount;                                    // F2H_Mem_Window_FF600000:avm_m0_burstcount -> mm_interconnect_1:F2H_Mem_Window_FF600000_expanded_master_burstcount
	wire         f2h_mem_window_ff800000_expanded_master_waitrequest;                                   // mm_interconnect_1:F2H_Mem_Window_FF800000_expanded_master_waitrequest -> F2H_Mem_Window_FF800000:avm_m0_waitrequest
	wire  [31:0] f2h_mem_window_ff800000_expanded_master_readdata;                                      // mm_interconnect_1:F2H_Mem_Window_FF800000_expanded_master_readdata -> F2H_Mem_Window_FF800000:avm_m0_readdata
	wire  [31:0] f2h_mem_window_ff800000_expanded_master_address;                                       // F2H_Mem_Window_FF800000:avm_m0_address -> mm_interconnect_1:F2H_Mem_Window_FF800000_expanded_master_address
	wire         f2h_mem_window_ff800000_expanded_master_read;                                          // F2H_Mem_Window_FF800000:avm_m0_read -> mm_interconnect_1:F2H_Mem_Window_FF800000_expanded_master_read
	wire   [3:0] f2h_mem_window_ff800000_expanded_master_byteenable;                                    // F2H_Mem_Window_FF800000:avm_m0_byteenable -> mm_interconnect_1:F2H_Mem_Window_FF800000_expanded_master_byteenable
	wire         f2h_mem_window_ff800000_expanded_master_readdatavalid;                                 // mm_interconnect_1:F2H_Mem_Window_FF800000_expanded_master_readdatavalid -> F2H_Mem_Window_FF800000:avm_m0_readdatavalid
	wire         f2h_mem_window_ff800000_expanded_master_write;                                         // F2H_Mem_Window_FF800000:avm_m0_write -> mm_interconnect_1:F2H_Mem_Window_FF800000_expanded_master_write
	wire  [31:0] f2h_mem_window_ff800000_expanded_master_writedata;                                     // F2H_Mem_Window_FF800000:avm_m0_writedata -> mm_interconnect_1:F2H_Mem_Window_FF800000_expanded_master_writedata
	wire   [0:0] f2h_mem_window_ff800000_expanded_master_burstcount;                                    // F2H_Mem_Window_FF800000:avm_m0_burstcount -> mm_interconnect_1:F2H_Mem_Window_FF800000_expanded_master_burstcount
	wire  [31:0] jtag_to_hps_bridge_master_readdata;                                                    // mm_interconnect_1:JTAG_to_HPS_Bridge_master_readdata -> JTAG_to_HPS_Bridge:master_readdata
	wire         jtag_to_hps_bridge_master_waitrequest;                                                 // mm_interconnect_1:JTAG_to_HPS_Bridge_master_waitrequest -> JTAG_to_HPS_Bridge:master_waitrequest
	wire  [31:0] jtag_to_hps_bridge_master_address;                                                     // JTAG_to_HPS_Bridge:master_address -> mm_interconnect_1:JTAG_to_HPS_Bridge_master_address
	wire         jtag_to_hps_bridge_master_read;                                                        // JTAG_to_HPS_Bridge:master_read -> mm_interconnect_1:JTAG_to_HPS_Bridge_master_read
	wire   [3:0] jtag_to_hps_bridge_master_byteenable;                                                  // JTAG_to_HPS_Bridge:master_byteenable -> mm_interconnect_1:JTAG_to_HPS_Bridge_master_byteenable
	wire         jtag_to_hps_bridge_master_readdatavalid;                                               // mm_interconnect_1:JTAG_to_HPS_Bridge_master_readdatavalid -> JTAG_to_HPS_Bridge:master_readdatavalid
	wire         jtag_to_hps_bridge_master_write;                                                       // JTAG_to_HPS_Bridge:master_write -> mm_interconnect_1:JTAG_to_HPS_Bridge_master_write
	wire  [31:0] jtag_to_hps_bridge_master_writedata;                                                   // JTAG_to_HPS_Bridge:master_writedata -> mm_interconnect_1:JTAG_to_HPS_Bridge_master_writedata
	wire   [1:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awburst;                                    // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awburst -> ARM_A9_HPS:f2h_AWBURST
	wire   [4:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awuser;                                     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awuser -> ARM_A9_HPS:f2h_AWUSER
	wire   [3:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlen;                                      // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arlen -> ARM_A9_HPS:f2h_ARLEN
	wire   [7:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wstrb;                                      // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wstrb -> ARM_A9_HPS:f2h_WSTRB
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wready;                                     // ARM_A9_HPS:f2h_WREADY -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wready
	wire   [7:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rid;                                        // ARM_A9_HPS:f2h_RID -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rid
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rready;                                     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rready -> ARM_A9_HPS:f2h_RREADY
	wire   [3:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlen;                                      // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awlen -> ARM_A9_HPS:f2h_AWLEN
	wire   [7:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wid;                                        // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wid -> ARM_A9_HPS:f2h_WID
	wire   [3:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arcache;                                    // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arcache -> ARM_A9_HPS:f2h_ARCACHE
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wvalid;                                     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wvalid -> ARM_A9_HPS:f2h_WVALID
	wire  [31:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_araddr;                                     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_araddr -> ARM_A9_HPS:f2h_ARADDR
	wire   [2:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arprot;                                     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arprot -> ARM_A9_HPS:f2h_ARPROT
	wire   [2:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awprot;                                     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awprot -> ARM_A9_HPS:f2h_AWPROT
	wire  [63:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wdata;                                      // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wdata -> ARM_A9_HPS:f2h_WDATA
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arvalid;                                    // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arvalid -> ARM_A9_HPS:f2h_ARVALID
	wire   [3:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awcache;                                    // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awcache -> ARM_A9_HPS:f2h_AWCACHE
	wire   [7:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arid;                                       // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arid -> ARM_A9_HPS:f2h_ARID
	wire   [1:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlock;                                     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arlock -> ARM_A9_HPS:f2h_ARLOCK
	wire   [1:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlock;                                     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awlock -> ARM_A9_HPS:f2h_AWLOCK
	wire  [31:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awaddr;                                     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awaddr -> ARM_A9_HPS:f2h_AWADDR
	wire   [1:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bresp;                                      // ARM_A9_HPS:f2h_BRESP -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_bresp
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arready;                                    // ARM_A9_HPS:f2h_ARREADY -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arready
	wire  [63:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rdata;                                      // ARM_A9_HPS:f2h_RDATA -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rdata
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awready;                                    // ARM_A9_HPS:f2h_AWREADY -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awready
	wire   [1:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arburst;                                    // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arburst -> ARM_A9_HPS:f2h_ARBURST
	wire   [2:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arsize;                                     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arsize -> ARM_A9_HPS:f2h_ARSIZE
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bready;                                     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_bready -> ARM_A9_HPS:f2h_BREADY
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rlast;                                      // ARM_A9_HPS:f2h_RLAST -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rlast
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wlast;                                      // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wlast -> ARM_A9_HPS:f2h_WLAST
	wire   [1:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rresp;                                      // ARM_A9_HPS:f2h_RRESP -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rresp
	wire   [7:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awid;                                       // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awid -> ARM_A9_HPS:f2h_AWID
	wire   [7:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bid;                                        // ARM_A9_HPS:f2h_BID -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_bid
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bvalid;                                     // ARM_A9_HPS:f2h_BVALID -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_bvalid
	wire   [2:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awsize;                                     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awsize -> ARM_A9_HPS:f2h_AWSIZE
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awvalid;                                    // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awvalid -> ARM_A9_HPS:f2h_AWVALID
	wire   [4:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_aruser;                                     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_aruser -> ARM_A9_HPS:f2h_ARUSER
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rvalid;                                     // ARM_A9_HPS:f2h_RVALID -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rvalid
	wire         irq_mapper_receiver6_irq;                                                              // JTAG_UART_for_ARM_0:av_irq -> irq_mapper:receiver6_irq
	wire  [31:0] arm_a9_hps_f2h_irq0_irq;                                                               // irq_mapper:sender_irq -> ARM_A9_HPS:f2h_irq_p0
	wire         irq_mapper_001_receiver0_irq;                                                          // JTAG_UART_for_ARM_1:av_irq -> irq_mapper_001:receiver0_irq
	wire  [31:0] arm_a9_hps_f2h_irq1_irq;                                                               // irq_mapper_001:sender_irq -> ARM_A9_HPS:f2h_irq_p1
	wire         irq_mapper_002_receiver6_irq;                                                          // JTAG_UART:av_irq -> irq_mapper_002:receiver6_irq
	wire  [31:0] nios2_irq_irq;                                                                         // irq_mapper_002:sender_irq -> Nios2:irq
	wire         irq_mapper_003_receiver6_irq;                                                          // JTAG_UART_2nd_Core:av_irq -> irq_mapper_003:receiver6_irq
	wire         irq_mapper_003_receiver7_irq;                                                          // Interval_Timer_2nd_Core:irq -> irq_mapper_003:receiver7_irq
	wire         irq_mapper_003_receiver8_irq;                                                          // Interval_Timer_2nd_Core_2:irq -> irq_mapper_003:receiver8_irq
	wire  [31:0] nios2_2nd_core_irq_irq;                                                                // irq_mapper_003:sender_irq -> Nios2_2nd_Core:irq
	wire         irq_mapper_receiver0_irq;                                                              // Audio_Subsystem:audio_irq_irq -> [irq_mapper:receiver0_irq, irq_mapper_002:receiver0_irq, irq_mapper_003:receiver0_irq]
	wire         irq_mapper_receiver5_irq;                                                              // Expansion_JP1:irq -> [irq_mapper:receiver5_irq, irq_mapper_002:receiver5_irq, irq_mapper_003:receiver5_irq]
	wire         irq_mapper_receiver7_irq;                                                              // Interval_Timer:irq -> [irq_mapper:receiver7_irq, irq_mapper_002:receiver7_irq]
	wire         irq_mapper_receiver8_irq;                                                              // Interval_Timer_2:irq -> [irq_mapper:receiver8_irq, irq_mapper_002:receiver8_irq]
	wire         irq_mapper_receiver3_irq;                                                              // IrDA:irq -> [irq_mapper:receiver3_irq, irq_mapper_002:receiver3_irq, irq_mapper_003:receiver3_irq]
	wire         irq_mapper_receiver1_irq;                                                              // PS2_Port:irq -> [irq_mapper:receiver1_irq, irq_mapper_002:receiver1_irq, irq_mapper_003:receiver1_irq]
	wire         irq_mapper_receiver2_irq;                                                              // PS2_Port_Dual:irq -> [irq_mapper:receiver2_irq, irq_mapper_002:receiver2_irq, irq_mapper_003:receiver2_irq]
	wire         irq_mapper_receiver4_irq;                                                              // Pushbuttons:irq -> [irq_mapper:receiver4_irq, irq_mapper_002:receiver4_irq, irq_mapper_003:receiver4_irq]
	wire         rst_controller_reset_out_reset;                                                        // rst_controller:reset_out -> [ADC:reset, AV_Config:reset, Char_DMA_Addr_Translation:reset, Expansion_JP1:reset_n, F2H_Mem_Window_00000000:reset, F2H_Mem_Window_FF600000:reset, F2H_Mem_Window_FF800000:reset, HEX3_HEX0:reset_n, HEX5_HEX4:reset_n, Interval_Timer:reset_n, Interval_Timer_2:reset_n, Interval_Timer_2nd_Core:reset_n, Interval_Timer_2nd_Core_2:reset_n, IrDA:reset, JTAG_UART:rst_n, JTAG_UART_2nd_Core:rst_n, JTAG_UART_for_ARM_0:rst_n, JTAG_UART_for_ARM_1:rst_n, LEDs:reset_n, Onchip_SRAM:reset, PS2_Port:reset, PS2_Port_Dual:reset, Pixel_DMA_Addr_Translation:reset, Pushbuttons:reset_n, SDRAM:reset_n, Slider_Switches:reset_n, SysID:reset_n, Video_In_DMA_Addr_Translation:reset, mm_interconnect_0:JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:Video_In_DMA_Addr_Translation_reset_reset_bridge_in_reset_reset, mm_interconnect_1:F2H_Mem_Window_00000000_reset_reset_bridge_in_reset_reset, mm_interconnect_1:JTAG_to_HPS_Bridge_clk_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                                                    // rst_controller:reset_req -> [Onchip_SRAM:reset_req, rst_translator:reset_req_in]
	wire         arm_a9_hps_h2f_reset_reset;                                                            // ARM_A9_HPS:h2f_rst_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0, rst_controller_004:reset_in1, rst_controller_005:reset_in1, rst_controller_006:reset_in0, rst_controller_007:reset_in0, rst_controller_008:reset_in0]
	wire         system_pll_reset_source_reset;                                                         // System_PLL:reset_source_reset -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1, rst_controller_004:reset_in2, rst_controller_005:reset_in2, rst_controller_006:reset_in1, rst_controller_007:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                                    // rst_controller_001:reset_out -> Audio_Subsystem:sys_reset_reset_n
	wire         rst_controller_002_reset_out_reset;                                                    // rst_controller_002:reset_out -> JTAG_to_FPGA_Bridge:clk_reset_reset
	wire         rst_controller_003_reset_out_reset;                                                    // rst_controller_003:reset_out -> JTAG_to_HPS_Bridge:clk_reset_reset
	wire         rst_controller_004_reset_out_reset;                                                    // rst_controller_004:reset_out -> [Nios2:reset_n, irq_mapper_002:reset, mm_interconnect_0:Nios2_reset_reset_bridge_in_reset_reset]
	wire         nios2_debug_reset_request_reset;                                                       // Nios2:debug_reset_request -> rst_controller_004:reset_in0
	wire         rst_controller_005_reset_out_reset;                                                    // rst_controller_005:reset_out -> [Nios2_2nd_Core:reset_n, irq_mapper_003:reset, mm_interconnect_0:Nios2_2nd_Core_reset_reset_bridge_in_reset_reset]
	wire         nios2_2nd_core_debug_reset_request_reset;                                              // Nios2_2nd_Core:debug_reset_request -> rst_controller_005:reset_in0
	wire         rst_controller_006_reset_out_reset;                                                    // rst_controller_006:reset_out -> VGA_Subsystem:sys_reset_reset_n
	wire         rst_controller_007_reset_out_reset;                                                    // rst_controller_007:reset_out -> Video_In_Subsystem:sys_reset_reset_n
	wire         rst_controller_008_reset_out_reset;                                                    // rst_controller_008:reset_out -> [mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset]

	Computer_System_ADC #(
		.board          ("DE10-Standard"),
		.board_rev      ("Autodetect"),
		.tsclk          (8),
		.numch          (7),
		.max10pllmultby (1),
		.max10plldivby  (1)
	) adc (
		.clock       (system_pll_sys_clk_clk),                      //                clk.clk
		.reset       (rst_controller_reset_out_reset),              //              reset.reset
		.write       (mm_interconnect_0_adc_adc_slave_write),       //          adc_slave.write
		.readdata    (mm_interconnect_0_adc_adc_slave_readdata),    //                   .readdata
		.writedata   (mm_interconnect_0_adc_adc_slave_writedata),   //                   .writedata
		.address     (mm_interconnect_0_adc_adc_slave_address),     //                   .address
		.waitrequest (mm_interconnect_0_adc_adc_slave_waitrequest), //                   .waitrequest
		.read        (mm_interconnect_0_adc_adc_slave_read),        //                   .read
		.adc_sclk    (adc_sclk),                                    // external_interface.export
		.adc_cs_n    (adc_cs_n),                                    //                   .export
		.adc_dout    (adc_dout),                                    //                   .export
		.adc_din     (adc_din)                                      //                   .export
	);

	Computer_System_ARM_A9_HPS #(
		.F2S_Width (2),
		.S2F_Width (2)
	) arm_a9_hps (
		.f2h_stm_hwevents         (),                                                   // f2h_stm_hw_events.stm_hwevents
		.mem_a                    (memory_mem_a),                                       //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                                      //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                                      //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                                    //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                     //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                                    //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                                   //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                                   //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                                    //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                                 //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                      //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                     //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                                   //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                     //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                                      //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                                   //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK),                    //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),                      //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),                      //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),                      //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),                      //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),                      //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),                      //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),                       //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL),                    //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL),                    //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK),                    //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),                      //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),                      //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),                      //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_io_hps_io_qspi_inst_IO0),                        //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_io_hps_io_qspi_inst_IO1),                        //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_io_hps_io_qspi_inst_IO2),                        //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_io_hps_io_qspi_inst_IO3),                        //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_io_hps_io_qspi_inst_SS0),                        //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_io_hps_io_qspi_inst_CLK),                        //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),                        //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),                         //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),                         //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),                        //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),                         //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),                         //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),                         //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),                         //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),                         //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),                         //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),                         //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),                         //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),                         //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),                         //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),                        //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),                        //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),                        //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),                        //                  .hps_io_usb1_inst_NXT
		.hps_io_spim0_inst_CLK    (hps_io_hps_io_spim0_inst_CLK),                       //                  .hps_io_spim0_inst_CLK
		.hps_io_spim0_inst_MOSI   (hps_io_hps_io_spim0_inst_MOSI),                      //                  .hps_io_spim0_inst_MOSI
		.hps_io_spim0_inst_MISO   (hps_io_hps_io_spim0_inst_MISO),                      //                  .hps_io_spim0_inst_MISO
		.hps_io_spim0_inst_SS0    (hps_io_hps_io_spim0_inst_SS0),                       //                  .hps_io_spim0_inst_SS0
		.hps_io_spim1_inst_CLK    (hps_io_hps_io_spim1_inst_CLK),                       //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_io_hps_io_spim1_inst_MOSI),                      //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_io_hps_io_spim1_inst_MISO),                      //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_io_hps_io_spim1_inst_SS0),                       //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),                        //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),                        //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),                        //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),                        //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),                        //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),                        //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_io_hps_io_gpio_inst_GPIO09),                     //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_io_hps_io_gpio_inst_GPIO35),                     //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO37  (hps_io_hps_io_gpio_inst_GPIO37),                     //                  .hps_io_gpio_inst_GPIO37
		.hps_io_gpio_inst_GPIO40  (hps_io_hps_io_gpio_inst_GPIO40),                     //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO41  (hps_io_hps_io_gpio_inst_GPIO41),                     //                  .hps_io_gpio_inst_GPIO41
		.hps_io_gpio_inst_GPIO44  (hps_io_hps_io_gpio_inst_GPIO44),                     //                  .hps_io_gpio_inst_GPIO44
		.hps_io_gpio_inst_GPIO48  (hps_io_hps_io_gpio_inst_GPIO48),                     //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_io_hps_io_gpio_inst_GPIO53),                     //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_io_hps_io_gpio_inst_GPIO54),                     //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_io_hps_io_gpio_inst_GPIO61),                     //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (arm_a9_hps_h2f_reset_reset),                         //         h2f_reset.reset_n
		.h2f_axi_clk              (system_pll_sys_clk_clk),                             //     h2f_axi_clock.clk
		.h2f_AWID                 (arm_a9_hps_h2f_axi_master_awid),                     //    h2f_axi_master.awid
		.h2f_AWADDR               (arm_a9_hps_h2f_axi_master_awaddr),                   //                  .awaddr
		.h2f_AWLEN                (arm_a9_hps_h2f_axi_master_awlen),                    //                  .awlen
		.h2f_AWSIZE               (arm_a9_hps_h2f_axi_master_awsize),                   //                  .awsize
		.h2f_AWBURST              (arm_a9_hps_h2f_axi_master_awburst),                  //                  .awburst
		.h2f_AWLOCK               (arm_a9_hps_h2f_axi_master_awlock),                   //                  .awlock
		.h2f_AWCACHE              (arm_a9_hps_h2f_axi_master_awcache),                  //                  .awcache
		.h2f_AWPROT               (arm_a9_hps_h2f_axi_master_awprot),                   //                  .awprot
		.h2f_AWVALID              (arm_a9_hps_h2f_axi_master_awvalid),                  //                  .awvalid
		.h2f_AWREADY              (arm_a9_hps_h2f_axi_master_awready),                  //                  .awready
		.h2f_WID                  (arm_a9_hps_h2f_axi_master_wid),                      //                  .wid
		.h2f_WDATA                (arm_a9_hps_h2f_axi_master_wdata),                    //                  .wdata
		.h2f_WSTRB                (arm_a9_hps_h2f_axi_master_wstrb),                    //                  .wstrb
		.h2f_WLAST                (arm_a9_hps_h2f_axi_master_wlast),                    //                  .wlast
		.h2f_WVALID               (arm_a9_hps_h2f_axi_master_wvalid),                   //                  .wvalid
		.h2f_WREADY               (arm_a9_hps_h2f_axi_master_wready),                   //                  .wready
		.h2f_BID                  (arm_a9_hps_h2f_axi_master_bid),                      //                  .bid
		.h2f_BRESP                (arm_a9_hps_h2f_axi_master_bresp),                    //                  .bresp
		.h2f_BVALID               (arm_a9_hps_h2f_axi_master_bvalid),                   //                  .bvalid
		.h2f_BREADY               (arm_a9_hps_h2f_axi_master_bready),                   //                  .bready
		.h2f_ARID                 (arm_a9_hps_h2f_axi_master_arid),                     //                  .arid
		.h2f_ARADDR               (arm_a9_hps_h2f_axi_master_araddr),                   //                  .araddr
		.h2f_ARLEN                (arm_a9_hps_h2f_axi_master_arlen),                    //                  .arlen
		.h2f_ARSIZE               (arm_a9_hps_h2f_axi_master_arsize),                   //                  .arsize
		.h2f_ARBURST              (arm_a9_hps_h2f_axi_master_arburst),                  //                  .arburst
		.h2f_ARLOCK               (arm_a9_hps_h2f_axi_master_arlock),                   //                  .arlock
		.h2f_ARCACHE              (arm_a9_hps_h2f_axi_master_arcache),                  //                  .arcache
		.h2f_ARPROT               (arm_a9_hps_h2f_axi_master_arprot),                   //                  .arprot
		.h2f_ARVALID              (arm_a9_hps_h2f_axi_master_arvalid),                  //                  .arvalid
		.h2f_ARREADY              (arm_a9_hps_h2f_axi_master_arready),                  //                  .arready
		.h2f_RID                  (arm_a9_hps_h2f_axi_master_rid),                      //                  .rid
		.h2f_RDATA                (arm_a9_hps_h2f_axi_master_rdata),                    //                  .rdata
		.h2f_RRESP                (arm_a9_hps_h2f_axi_master_rresp),                    //                  .rresp
		.h2f_RLAST                (arm_a9_hps_h2f_axi_master_rlast),                    //                  .rlast
		.h2f_RVALID               (arm_a9_hps_h2f_axi_master_rvalid),                   //                  .rvalid
		.h2f_RREADY               (arm_a9_hps_h2f_axi_master_rready),                   //                  .rready
		.f2h_axi_clk              (system_pll_sys_clk_clk),                             //     f2h_axi_clock.clk
		.f2h_AWID                 (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awid),    //     f2h_axi_slave.awid
		.f2h_AWADDR               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awaddr),  //                  .awaddr
		.f2h_AWLEN                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlen),   //                  .awlen
		.f2h_AWSIZE               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awsize),  //                  .awsize
		.f2h_AWBURST              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awburst), //                  .awburst
		.f2h_AWLOCK               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlock),  //                  .awlock
		.f2h_AWCACHE              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awcache), //                  .awcache
		.f2h_AWPROT               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awprot),  //                  .awprot
		.f2h_AWVALID              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awvalid), //                  .awvalid
		.f2h_AWREADY              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awready), //                  .awready
		.f2h_AWUSER               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awuser),  //                  .awuser
		.f2h_WID                  (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wid),     //                  .wid
		.f2h_WDATA                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wdata),   //                  .wdata
		.f2h_WSTRB                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wstrb),   //                  .wstrb
		.f2h_WLAST                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wlast),   //                  .wlast
		.f2h_WVALID               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wvalid),  //                  .wvalid
		.f2h_WREADY               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wready),  //                  .wready
		.f2h_BID                  (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bid),     //                  .bid
		.f2h_BRESP                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bresp),   //                  .bresp
		.f2h_BVALID               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bvalid),  //                  .bvalid
		.f2h_BREADY               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bready),  //                  .bready
		.f2h_ARID                 (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arid),    //                  .arid
		.f2h_ARADDR               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_araddr),  //                  .araddr
		.f2h_ARLEN                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlen),   //                  .arlen
		.f2h_ARSIZE               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arsize),  //                  .arsize
		.f2h_ARBURST              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arburst), //                  .arburst
		.f2h_ARLOCK               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlock),  //                  .arlock
		.f2h_ARCACHE              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arcache), //                  .arcache
		.f2h_ARPROT               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arprot),  //                  .arprot
		.f2h_ARVALID              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arvalid), //                  .arvalid
		.f2h_ARREADY              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arready), //                  .arready
		.f2h_ARUSER               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_aruser),  //                  .aruser
		.f2h_RID                  (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rid),     //                  .rid
		.f2h_RDATA                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rdata),   //                  .rdata
		.f2h_RRESP                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rresp),   //                  .rresp
		.f2h_RLAST                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rlast),   //                  .rlast
		.f2h_RVALID               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rvalid),  //                  .rvalid
		.f2h_RREADY               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rready),  //                  .rready
		.h2f_lw_axi_clk           (system_pll_sys_clk_clk),                             //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (arm_a9_hps_h2f_lw_axi_master_awid),                  // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (arm_a9_hps_h2f_lw_axi_master_awaddr),                //                  .awaddr
		.h2f_lw_AWLEN             (arm_a9_hps_h2f_lw_axi_master_awlen),                 //                  .awlen
		.h2f_lw_AWSIZE            (arm_a9_hps_h2f_lw_axi_master_awsize),                //                  .awsize
		.h2f_lw_AWBURST           (arm_a9_hps_h2f_lw_axi_master_awburst),               //                  .awburst
		.h2f_lw_AWLOCK            (arm_a9_hps_h2f_lw_axi_master_awlock),                //                  .awlock
		.h2f_lw_AWCACHE           (arm_a9_hps_h2f_lw_axi_master_awcache),               //                  .awcache
		.h2f_lw_AWPROT            (arm_a9_hps_h2f_lw_axi_master_awprot),                //                  .awprot
		.h2f_lw_AWVALID           (arm_a9_hps_h2f_lw_axi_master_awvalid),               //                  .awvalid
		.h2f_lw_AWREADY           (arm_a9_hps_h2f_lw_axi_master_awready),               //                  .awready
		.h2f_lw_WID               (arm_a9_hps_h2f_lw_axi_master_wid),                   //                  .wid
		.h2f_lw_WDATA             (arm_a9_hps_h2f_lw_axi_master_wdata),                 //                  .wdata
		.h2f_lw_WSTRB             (arm_a9_hps_h2f_lw_axi_master_wstrb),                 //                  .wstrb
		.h2f_lw_WLAST             (arm_a9_hps_h2f_lw_axi_master_wlast),                 //                  .wlast
		.h2f_lw_WVALID            (arm_a9_hps_h2f_lw_axi_master_wvalid),                //                  .wvalid
		.h2f_lw_WREADY            (arm_a9_hps_h2f_lw_axi_master_wready),                //                  .wready
		.h2f_lw_BID               (arm_a9_hps_h2f_lw_axi_master_bid),                   //                  .bid
		.h2f_lw_BRESP             (arm_a9_hps_h2f_lw_axi_master_bresp),                 //                  .bresp
		.h2f_lw_BVALID            (arm_a9_hps_h2f_lw_axi_master_bvalid),                //                  .bvalid
		.h2f_lw_BREADY            (arm_a9_hps_h2f_lw_axi_master_bready),                //                  .bready
		.h2f_lw_ARID              (arm_a9_hps_h2f_lw_axi_master_arid),                  //                  .arid
		.h2f_lw_ARADDR            (arm_a9_hps_h2f_lw_axi_master_araddr),                //                  .araddr
		.h2f_lw_ARLEN             (arm_a9_hps_h2f_lw_axi_master_arlen),                 //                  .arlen
		.h2f_lw_ARSIZE            (arm_a9_hps_h2f_lw_axi_master_arsize),                //                  .arsize
		.h2f_lw_ARBURST           (arm_a9_hps_h2f_lw_axi_master_arburst),               //                  .arburst
		.h2f_lw_ARLOCK            (arm_a9_hps_h2f_lw_axi_master_arlock),                //                  .arlock
		.h2f_lw_ARCACHE           (arm_a9_hps_h2f_lw_axi_master_arcache),               //                  .arcache
		.h2f_lw_ARPROT            (arm_a9_hps_h2f_lw_axi_master_arprot),                //                  .arprot
		.h2f_lw_ARVALID           (arm_a9_hps_h2f_lw_axi_master_arvalid),               //                  .arvalid
		.h2f_lw_ARREADY           (arm_a9_hps_h2f_lw_axi_master_arready),               //                  .arready
		.h2f_lw_RID               (arm_a9_hps_h2f_lw_axi_master_rid),                   //                  .rid
		.h2f_lw_RDATA             (arm_a9_hps_h2f_lw_axi_master_rdata),                 //                  .rdata
		.h2f_lw_RRESP             (arm_a9_hps_h2f_lw_axi_master_rresp),                 //                  .rresp
		.h2f_lw_RLAST             (arm_a9_hps_h2f_lw_axi_master_rlast),                 //                  .rlast
		.h2f_lw_RVALID            (arm_a9_hps_h2f_lw_axi_master_rvalid),                //                  .rvalid
		.h2f_lw_RREADY            (arm_a9_hps_h2f_lw_axi_master_rready),                //                  .rready
		.f2h_irq_p0               (arm_a9_hps_f2h_irq0_irq),                            //          f2h_irq0.irq
		.f2h_irq_p1               (arm_a9_hps_f2h_irq1_irq)                             //          f2h_irq1.irq
	);

	Computer_System_AV_Config av_config (
		.clk         (system_pll_sys_clk_clk),                                         //                    clk.clk
		.reset       (rst_controller_reset_out_reset),                                 //                  reset.reset
		.address     (mm_interconnect_0_av_config_avalon_av_config_slave_address),     // avalon_av_config_slave.address
		.byteenable  (mm_interconnect_0_av_config_avalon_av_config_slave_byteenable),  //                       .byteenable
		.read        (mm_interconnect_0_av_config_avalon_av_config_slave_read),        //                       .read
		.write       (mm_interconnect_0_av_config_avalon_av_config_slave_write),       //                       .write
		.writedata   (mm_interconnect_0_av_config_avalon_av_config_slave_writedata),   //                       .writedata
		.readdata    (mm_interconnect_0_av_config_avalon_av_config_slave_readdata),    //                       .readdata
		.waitrequest (mm_interconnect_0_av_config_avalon_av_config_slave_waitrequest), //                       .waitrequest
		.I2C_SDAT    (av_config_SDAT),                                                 //     external_interface.export
		.I2C_SCLK    (av_config_SCLK)                                                  //                       .export
	);

	Computer_System_Audio_Subsystem audio_subsystem (
		.audio_ADCDAT              (audio_ADCDAT),                                             //               audio.ADCDAT
		.audio_ADCLRCK             (audio_ADCLRCK),                                            //                    .ADCLRCK
		.audio_BCLK                (audio_BCLK),                                               //                    .BCLK
		.audio_DACDAT              (audio_DACDAT),                                             //                    .DACDAT
		.audio_DACLRCK             (audio_DACLRCK),                                            //                    .DACLRCK
		.audio_irq_irq             (irq_mapper_receiver0_irq),                                 //           audio_irq.irq
		.audio_pll_clk_clk         (audio_pll_clk_clk),                                        //       audio_pll_clk.clk
		.audio_pll_ref_clk_clk     (audio_pll_ref_clk_clk),                                    //   audio_pll_ref_clk.clk
		.audio_pll_ref_reset_reset (audio_pll_ref_reset_reset),                                // audio_pll_ref_reset.reset
		.audio_pll_reset_reset     (),                                                         //     audio_pll_reset.reset
		.audio_slave_address       (mm_interconnect_0_audio_subsystem_audio_slave_address),    //         audio_slave.address
		.audio_slave_chipselect    (mm_interconnect_0_audio_subsystem_audio_slave_chipselect), //                    .chipselect
		.audio_slave_read          (mm_interconnect_0_audio_subsystem_audio_slave_read),       //                    .read
		.audio_slave_write         (mm_interconnect_0_audio_subsystem_audio_slave_write),      //                    .write
		.audio_slave_writedata     (mm_interconnect_0_audio_subsystem_audio_slave_writedata),  //                    .writedata
		.audio_slave_readdata      (mm_interconnect_0_audio_subsystem_audio_slave_readdata),   //                    .readdata
		.sys_clk_clk               (system_pll_sys_clk_clk),                                   //             sys_clk.clk
		.sys_reset_reset_n         (~rst_controller_001_reset_out_reset)                       //           sys_reset.reset_n
	);

	altera_up_avalon_video_dma_ctrl_addr_trans #(
		.ADDRESS_TRANSLATION_MASK (32'b11000000000000000000000000000000)
	) char_dma_addr_translation (
		.clk                (system_pll_sys_clk_clk),                                        //  clock.clk
		.reset              (rst_controller_reset_out_reset),                                //  reset.reset
		.slave_address      (mm_interconnect_0_char_dma_addr_translation_slave_address),     //  slave.address
		.slave_byteenable   (mm_interconnect_0_char_dma_addr_translation_slave_byteenable),  //       .byteenable
		.slave_read         (mm_interconnect_0_char_dma_addr_translation_slave_read),        //       .read
		.slave_write        (mm_interconnect_0_char_dma_addr_translation_slave_write),       //       .write
		.slave_writedata    (mm_interconnect_0_char_dma_addr_translation_slave_writedata),   //       .writedata
		.slave_readdata     (mm_interconnect_0_char_dma_addr_translation_slave_readdata),    //       .readdata
		.slave_waitrequest  (mm_interconnect_0_char_dma_addr_translation_slave_waitrequest), //       .waitrequest
		.master_readdata    (char_dma_addr_translation_master_readdata),                     // master.readdata
		.master_waitrequest (char_dma_addr_translation_master_waitrequest),                  //       .waitrequest
		.master_address     (char_dma_addr_translation_master_address),                      //       .address
		.master_byteenable  (char_dma_addr_translation_master_byteenable),                   //       .byteenable
		.master_read        (char_dma_addr_translation_master_read),                         //       .read
		.master_write       (char_dma_addr_translation_master_write),                        //       .write
		.master_writedata   (char_dma_addr_translation_master_writedata)                     //       .writedata
	);

	Computer_System_Expansion_JP1 expansion_jp1 (
		.clk        (system_pll_sys_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_expansion_jp1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_expansion_jp1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_expansion_jp1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_expansion_jp1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_expansion_jp1_s1_readdata),   //                    .readdata
		.bidir_port (expansion_jp1_export),                          // external_connection.export
		.irq        (irq_mapper_receiver5_irq)                       //                 irq.irq
	);

	altera_address_span_extender #(
		.DATA_WIDTH           (32),
		.BYTEENABLE_WIDTH     (4),
		.MASTER_ADDRESS_WIDTH (32),
		.SLAVE_ADDRESS_WIDTH  (28),
		.SLAVE_ADDRESS_SHIFT  (2),
		.BURSTCOUNT_WIDTH     (1),
		.CNTL_ADDRESS_WIDTH   (1),
		.SUB_WINDOW_COUNT     (1),
		.MASTER_ADDRESS_DEF   (64'b0000000000000000000000000000000000000000000000000000000000000000)
	) f2h_mem_window_00000000 (
		.clk                  (system_pll_sys_clk_clk),                                                 //           clock.clk
		.reset                (rst_controller_reset_out_reset),                                         //           reset.reset
		.avs_s0_address       (mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_address),       //  windowed_slave.address
		.avs_s0_read          (mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_read),          //                .read
		.avs_s0_readdata      (mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_readdata),      //                .readdata
		.avs_s0_write         (mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_write),         //                .write
		.avs_s0_writedata     (mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_writedata),     //                .writedata
		.avs_s0_readdatavalid (mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_readdatavalid), //                .readdatavalid
		.avs_s0_waitrequest   (mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_waitrequest),   //                .waitrequest
		.avs_s0_byteenable    (mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_byteenable),    //                .byteenable
		.avs_s0_burstcount    (mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_burstcount),    //                .burstcount
		.avm_m0_address       (f2h_mem_window_00000000_expanded_master_address),                        // expanded_master.address
		.avm_m0_read          (f2h_mem_window_00000000_expanded_master_read),                           //                .read
		.avm_m0_waitrequest   (f2h_mem_window_00000000_expanded_master_waitrequest),                    //                .waitrequest
		.avm_m0_readdata      (f2h_mem_window_00000000_expanded_master_readdata),                       //                .readdata
		.avm_m0_write         (f2h_mem_window_00000000_expanded_master_write),                          //                .write
		.avm_m0_writedata     (f2h_mem_window_00000000_expanded_master_writedata),                      //                .writedata
		.avm_m0_readdatavalid (f2h_mem_window_00000000_expanded_master_readdatavalid),                  //                .readdatavalid
		.avm_m0_byteenable    (f2h_mem_window_00000000_expanded_master_byteenable),                     //                .byteenable
		.avm_m0_burstcount    (f2h_mem_window_00000000_expanded_master_burstcount),                     //                .burstcount
		.avs_cntl_address     (1'b0),                                                                   //     (terminated)
		.avs_cntl_read        (1'b0),                                                                   //     (terminated)
		.avs_cntl_readdata    (),                                                                       //     (terminated)
		.avs_cntl_write       (1'b0),                                                                   //     (terminated)
		.avs_cntl_writedata   (64'b0000000000000000000000000000000000000000000000000000000000000000),   //     (terminated)
		.avs_cntl_byteenable  (8'b00000000)                                                             //     (terminated)
	);

	altera_address_span_extender #(
		.DATA_WIDTH           (32),
		.BYTEENABLE_WIDTH     (4),
		.MASTER_ADDRESS_WIDTH (32),
		.SLAVE_ADDRESS_WIDTH  (19),
		.SLAVE_ADDRESS_SHIFT  (2),
		.BURSTCOUNT_WIDTH     (1),
		.CNTL_ADDRESS_WIDTH   (1),
		.SUB_WINDOW_COUNT     (1),
		.MASTER_ADDRESS_DEF   (64'b0000000000000000000000000000000011111111011000000000000000000000)
	) f2h_mem_window_ff600000 (
		.clk                  (system_pll_sys_clk_clk),                                                 //           clock.clk
		.reset                (rst_controller_reset_out_reset),                                         //           reset.reset
		.avs_s0_address       (mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_address),       //  windowed_slave.address
		.avs_s0_read          (mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_read),          //                .read
		.avs_s0_readdata      (mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_readdata),      //                .readdata
		.avs_s0_write         (mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_write),         //                .write
		.avs_s0_writedata     (mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_writedata),     //                .writedata
		.avs_s0_readdatavalid (mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_readdatavalid), //                .readdatavalid
		.avs_s0_waitrequest   (mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_waitrequest),   //                .waitrequest
		.avs_s0_byteenable    (mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_byteenable),    //                .byteenable
		.avs_s0_burstcount    (mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_burstcount),    //                .burstcount
		.avm_m0_address       (f2h_mem_window_ff600000_expanded_master_address),                        // expanded_master.address
		.avm_m0_read          (f2h_mem_window_ff600000_expanded_master_read),                           //                .read
		.avm_m0_waitrequest   (f2h_mem_window_ff600000_expanded_master_waitrequest),                    //                .waitrequest
		.avm_m0_readdata      (f2h_mem_window_ff600000_expanded_master_readdata),                       //                .readdata
		.avm_m0_write         (f2h_mem_window_ff600000_expanded_master_write),                          //                .write
		.avm_m0_writedata     (f2h_mem_window_ff600000_expanded_master_writedata),                      //                .writedata
		.avm_m0_readdatavalid (f2h_mem_window_ff600000_expanded_master_readdatavalid),                  //                .readdatavalid
		.avm_m0_byteenable    (f2h_mem_window_ff600000_expanded_master_byteenable),                     //                .byteenable
		.avm_m0_burstcount    (f2h_mem_window_ff600000_expanded_master_burstcount),                     //                .burstcount
		.avs_cntl_address     (1'b0),                                                                   //     (terminated)
		.avs_cntl_read        (1'b0),                                                                   //     (terminated)
		.avs_cntl_readdata    (),                                                                       //     (terminated)
		.avs_cntl_write       (1'b0),                                                                   //     (terminated)
		.avs_cntl_writedata   (64'b0000000000000000000000000000000000000000000000000000000000000000),   //     (terminated)
		.avs_cntl_byteenable  (8'b00000000)                                                             //     (terminated)
	);

	altera_address_span_extender #(
		.DATA_WIDTH           (32),
		.BYTEENABLE_WIDTH     (4),
		.MASTER_ADDRESS_WIDTH (32),
		.SLAVE_ADDRESS_WIDTH  (21),
		.SLAVE_ADDRESS_SHIFT  (2),
		.BURSTCOUNT_WIDTH     (1),
		.CNTL_ADDRESS_WIDTH   (1),
		.SUB_WINDOW_COUNT     (1),
		.MASTER_ADDRESS_DEF   (64'b0000000000000000000000000000000011111111100000000000000000000000)
	) f2h_mem_window_ff800000 (
		.clk                  (system_pll_sys_clk_clk),                                                 //           clock.clk
		.reset                (rst_controller_reset_out_reset),                                         //           reset.reset
		.avs_s0_address       (mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_address),       //  windowed_slave.address
		.avs_s0_read          (mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_read),          //                .read
		.avs_s0_readdata      (mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_readdata),      //                .readdata
		.avs_s0_write         (mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_write),         //                .write
		.avs_s0_writedata     (mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_writedata),     //                .writedata
		.avs_s0_readdatavalid (mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_readdatavalid), //                .readdatavalid
		.avs_s0_waitrequest   (mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_waitrequest),   //                .waitrequest
		.avs_s0_byteenable    (mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_byteenable),    //                .byteenable
		.avs_s0_burstcount    (mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_burstcount),    //                .burstcount
		.avm_m0_address       (f2h_mem_window_ff800000_expanded_master_address),                        // expanded_master.address
		.avm_m0_read          (f2h_mem_window_ff800000_expanded_master_read),                           //                .read
		.avm_m0_waitrequest   (f2h_mem_window_ff800000_expanded_master_waitrequest),                    //                .waitrequest
		.avm_m0_readdata      (f2h_mem_window_ff800000_expanded_master_readdata),                       //                .readdata
		.avm_m0_write         (f2h_mem_window_ff800000_expanded_master_write),                          //                .write
		.avm_m0_writedata     (f2h_mem_window_ff800000_expanded_master_writedata),                      //                .writedata
		.avm_m0_readdatavalid (f2h_mem_window_ff800000_expanded_master_readdatavalid),                  //                .readdatavalid
		.avm_m0_byteenable    (f2h_mem_window_ff800000_expanded_master_byteenable),                     //                .byteenable
		.avm_m0_burstcount    (f2h_mem_window_ff800000_expanded_master_burstcount),                     //                .burstcount
		.avs_cntl_address     (1'b0),                                                                   //     (terminated)
		.avs_cntl_read        (1'b0),                                                                   //     (terminated)
		.avs_cntl_readdata    (),                                                                       //     (terminated)
		.avs_cntl_write       (1'b0),                                                                   //     (terminated)
		.avs_cntl_writedata   (64'b0000000000000000000000000000000000000000000000000000000000000000),   //     (terminated)
		.avs_cntl_byteenable  (8'b00000000)                                                             //     (terminated)
	);

	Computer_System_HEX3_HEX0 hex3_hex0 (
		.clk        (system_pll_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_hex3_hex0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex3_hex0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex3_hex0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex3_hex0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex3_hex0_s1_readdata),   //                    .readdata
		.out_port   (hex3_hex0_export)                           // external_connection.export
	);

	Computer_System_HEX5_HEX4 hex5_hex4 (
		.clk        (system_pll_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_hex5_hex4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex5_hex4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex5_hex4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex5_hex4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex5_hex4_s1_readdata),   //                    .readdata
		.out_port   (hex5_hex4_export)                           // external_connection.export
	);

	Computer_System_Interval_Timer interval_timer (
		.clk        (system_pll_sys_clk_clk),                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                // reset.reset_n
		.address    (mm_interconnect_0_interval_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_interval_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_interval_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_interval_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_interval_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver7_irq)                        //   irq.irq
	);

	Computer_System_Interval_Timer interval_timer_2 (
		.clk        (system_pll_sys_clk_clk),                           //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  // reset.reset_n
		.address    (mm_interconnect_0_interval_timer_2_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_interval_timer_2_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_interval_timer_2_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_interval_timer_2_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_interval_timer_2_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver8_irq)                          //   irq.irq
	);

	Computer_System_Interval_Timer interval_timer_2nd_core (
		.clk        (system_pll_sys_clk_clk),                                  //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                         // reset.reset_n
		.address    (mm_interconnect_0_interval_timer_2nd_core_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_interval_timer_2nd_core_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_interval_timer_2nd_core_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_interval_timer_2nd_core_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_interval_timer_2nd_core_s1_write),     //      .write_n
		.irq        (irq_mapper_003_receiver7_irq)                             //   irq.irq
	);

	Computer_System_Interval_Timer interval_timer_2nd_core_2 (
		.clk        (system_pll_sys_clk_clk),                                    //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                           // reset.reset_n
		.address    (mm_interconnect_0_interval_timer_2nd_core_2_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_interval_timer_2nd_core_2_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_interval_timer_2nd_core_2_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_interval_timer_2nd_core_2_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_interval_timer_2nd_core_2_s1_write),     //      .write_n
		.irq        (irq_mapper_003_receiver8_irq)                               //   irq.irq
	);

	Computer_System_IrDA irda (
		.clk        (system_pll_sys_clk_clk),                              //                clk.clk
		.reset      (rst_controller_reset_out_reset),                      //              reset.reset
		.address    (mm_interconnect_0_irda_avalon_irda_slave_address),    //  avalon_irda_slave.address
		.chipselect (mm_interconnect_0_irda_avalon_irda_slave_chipselect), //                   .chipselect
		.byteenable (mm_interconnect_0_irda_avalon_irda_slave_byteenable), //                   .byteenable
		.read       (mm_interconnect_0_irda_avalon_irda_slave_read),       //                   .read
		.write      (mm_interconnect_0_irda_avalon_irda_slave_write),      //                   .write
		.writedata  (mm_interconnect_0_irda_avalon_irda_slave_writedata),  //                   .writedata
		.readdata   (mm_interconnect_0_irda_avalon_irda_slave_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver3_irq),                            //          interrupt.irq
		.IRDA_TXD   (irda_TXD),                                            // external_interface.export
		.IRDA_RXD   (irda_RXD)                                             //                   .export
	);

	Computer_System_JTAG_UART jtag_uart (
		.clk            (system_pll_sys_clk_clk),                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_002_receiver6_irq)                               //               irq.irq
	);

	Computer_System_JTAG_UART jtag_uart_2nd_core (
		.clk            (system_pll_sys_clk_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                    //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_003_receiver6_irq)                                        //               irq.irq
	);

	Computer_System_JTAG_UART jtag_uart_for_arm_0 (
		.clk            (system_pll_sys_clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                     //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver6_irq)                                             //               irq.irq
	);

	Computer_System_JTAG_UART jtag_uart_for_arm_1 (
		.clk            (system_pll_sys_clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                     //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver0_irq)                                         //               irq.irq
	);

	Computer_System_JTAG_to_FPGA_Bridge #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) jtag_to_fpga_bridge (
		.clk_clk              (system_pll_sys_clk_clk),                   //          clk.clk
		.clk_reset_reset      (rst_controller_002_reset_out_reset),       //    clk_reset.reset
		.master_address       (jtag_to_fpga_bridge_master_address),       //       master.address
		.master_readdata      (jtag_to_fpga_bridge_master_readdata),      //             .readdata
		.master_read          (jtag_to_fpga_bridge_master_read),          //             .read
		.master_write         (jtag_to_fpga_bridge_master_write),         //             .write
		.master_writedata     (jtag_to_fpga_bridge_master_writedata),     //             .writedata
		.master_waitrequest   (jtag_to_fpga_bridge_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (jtag_to_fpga_bridge_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (jtag_to_fpga_bridge_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                          // master_reset.reset
	);

	Computer_System_JTAG_to_FPGA_Bridge #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) jtag_to_hps_bridge (
		.clk_clk              (system_pll_sys_clk_clk),                  //          clk.clk
		.clk_reset_reset      (rst_controller_003_reset_out_reset),      //    clk_reset.reset
		.master_address       (jtag_to_hps_bridge_master_address),       //       master.address
		.master_readdata      (jtag_to_hps_bridge_master_readdata),      //             .readdata
		.master_read          (jtag_to_hps_bridge_master_read),          //             .read
		.master_write         (jtag_to_hps_bridge_master_write),         //             .write
		.master_writedata     (jtag_to_hps_bridge_master_writedata),     //             .writedata
		.master_waitrequest   (jtag_to_hps_bridge_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (jtag_to_hps_bridge_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (jtag_to_hps_bridge_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                         // master_reset.reset
	);

	Computer_System_LEDs leds (
		.clk        (system_pll_sys_clk_clk),               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	Computer_System_Nios2 nios2 (
		.clk                                 (system_pll_sys_clk_clk),                              //                       clk.clk
		.reset_n                             (~rst_controller_004_reset_out_reset),                 //                     reset.reset_n
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.A_ci_multi_done                     (nios2_custom_instruction_master_done),                // custom_instruction_master.done
		.A_ci_multi_result                   (nios2_custom_instruction_master_multi_result),        //                          .multi_result
		.A_ci_multi_a                        (nios2_custom_instruction_master_multi_a),             //                          .multi_a
		.A_ci_multi_b                        (nios2_custom_instruction_master_multi_b),             //                          .multi_b
		.A_ci_multi_c                        (nios2_custom_instruction_master_multi_c),             //                          .multi_c
		.A_ci_multi_clk_en                   (nios2_custom_instruction_master_clk_en),              //                          .clk_en
		.A_ci_multi_clock                    (nios2_custom_instruction_master_clk),                 //                          .clk
		.A_ci_multi_reset                    (nios2_custom_instruction_master_reset),               //                          .reset
		.A_ci_multi_reset_req                (nios2_custom_instruction_master_reset_req),           //                          .reset_req
		.A_ci_multi_dataa                    (nios2_custom_instruction_master_multi_dataa),         //                          .multi_dataa
		.A_ci_multi_datab                    (nios2_custom_instruction_master_multi_datab),         //                          .multi_datab
		.A_ci_multi_n                        (nios2_custom_instruction_master_multi_n),             //                          .multi_n
		.A_ci_multi_readra                   (nios2_custom_instruction_master_multi_readra),        //                          .multi_readra
		.A_ci_multi_readrb                   (nios2_custom_instruction_master_multi_readrb),        //                          .multi_readrb
		.A_ci_multi_start                    (nios2_custom_instruction_master_start),               //                          .start
		.A_ci_multi_writerc                  (nios2_custom_instruction_master_multi_writerc)        //                          .multi_writerc
	);

	Computer_System_Nios2_2nd_Core nios2_2nd_core (
		.clk                                 (system_pll_sys_clk_clk),                                       //                       clk.clk
		.reset_n                             (~rst_controller_005_reset_out_reset),                          //                     reset.reset_n
		.d_address                           (nios2_2nd_core_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_2nd_core_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_2nd_core_data_master_read),                              //                          .read
		.d_readdata                          (nios2_2nd_core_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_2nd_core_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_2nd_core_data_master_write),                             //                          .write
		.d_writedata                         (nios2_2nd_core_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_2nd_core_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_2nd_core_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_2nd_core_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_2nd_core_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_2nd_core_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_2nd_core_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_2nd_core_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_2nd_core_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_writedata),   //                          .writedata
		.A_ci_multi_done                     (nios2_2nd_core_custom_instruction_master_done),                // custom_instruction_master.done
		.A_ci_multi_result                   (nios2_2nd_core_custom_instruction_master_multi_result),        //                          .multi_result
		.A_ci_multi_a                        (nios2_2nd_core_custom_instruction_master_multi_a),             //                          .multi_a
		.A_ci_multi_b                        (nios2_2nd_core_custom_instruction_master_multi_b),             //                          .multi_b
		.A_ci_multi_c                        (nios2_2nd_core_custom_instruction_master_multi_c),             //                          .multi_c
		.A_ci_multi_clk_en                   (nios2_2nd_core_custom_instruction_master_clk_en),              //                          .clk_en
		.A_ci_multi_clock                    (nios2_2nd_core_custom_instruction_master_clk),                 //                          .clk
		.A_ci_multi_reset                    (nios2_2nd_core_custom_instruction_master_reset),               //                          .reset
		.A_ci_multi_reset_req                (nios2_2nd_core_custom_instruction_master_reset_req),           //                          .reset_req
		.A_ci_multi_dataa                    (nios2_2nd_core_custom_instruction_master_multi_dataa),         //                          .multi_dataa
		.A_ci_multi_datab                    (nios2_2nd_core_custom_instruction_master_multi_datab),         //                          .multi_datab
		.A_ci_multi_n                        (nios2_2nd_core_custom_instruction_master_multi_n),             //                          .multi_n
		.A_ci_multi_readra                   (nios2_2nd_core_custom_instruction_master_multi_readra),        //                          .multi_readra
		.A_ci_multi_readrb                   (nios2_2nd_core_custom_instruction_master_multi_readrb),        //                          .multi_readrb
		.A_ci_multi_start                    (nios2_2nd_core_custom_instruction_master_start),               //                          .start
		.A_ci_multi_writerc                  (nios2_2nd_core_custom_instruction_master_multi_writerc)        //                          .multi_writerc
	);

	fpoint_wrapper #(
		.useDivider (1)
	) nios2_2nd_core_floating_point (
		.clk    (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_clk),    // s1.clk
		.clk_en (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //   .clk_en
		.dataa  (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  //   .dataa
		.datab  (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //   .datab
		.n      (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_n),      //   .n
		.reset  (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //   .reset
		.start  (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_start),  //   .start
		.done   (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_done),   //   .done
		.result (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_result)  //   .result
	);

	fpoint_wrapper #(
		.useDivider (1)
	) nios2_floating_point (
		.clk    (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk),    // s1.clk
		.clk_en (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //   .clk_en
		.dataa  (nios2_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  //   .dataa
		.datab  (nios2_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //   .datab
		.n      (nios2_custom_instruction_master_multi_slave_translator0_ci_master_n),      //   .n
		.reset  (nios2_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //   .reset
		.start  (nios2_custom_instruction_master_multi_slave_translator0_ci_master_start),  //   .start
		.done   (nios2_custom_instruction_master_multi_slave_translator0_ci_master_done),   //   .done
		.result (nios2_custom_instruction_master_multi_slave_translator0_ci_master_result)  //   .result
	);

	Computer_System_Onchip_SRAM onchip_sram (
		.address     (mm_interconnect_0_onchip_sram_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_onchip_sram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_onchip_sram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_onchip_sram_s1_write),      //       .write
		.readdata    (mm_interconnect_0_onchip_sram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_onchip_sram_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_onchip_sram_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_0_onchip_sram_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_onchip_sram_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_onchip_sram_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_onchip_sram_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_onchip_sram_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_onchip_sram_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_onchip_sram_s2_byteenable), //       .byteenable
		.clk         (system_pll_sys_clk_clk),                      //   clk1.clk
		.reset       (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),          //       .reset_req
		.freeze      (1'b0)                                         // (terminated)
	);

	Computer_System_PS2_Port ps2_port (
		.clk         (system_pll_sys_clk_clk),                                  //                clk.clk
		.reset       (rst_controller_reset_out_reset),                          //              reset.reset
		.address     (mm_interconnect_0_ps2_port_avalon_ps2_slave_address),     //   avalon_ps2_slave.address
		.chipselect  (mm_interconnect_0_ps2_port_avalon_ps2_slave_chipselect),  //                   .chipselect
		.byteenable  (mm_interconnect_0_ps2_port_avalon_ps2_slave_byteenable),  //                   .byteenable
		.read        (mm_interconnect_0_ps2_port_avalon_ps2_slave_read),        //                   .read
		.write       (mm_interconnect_0_ps2_port_avalon_ps2_slave_write),       //                   .write
		.writedata   (mm_interconnect_0_ps2_port_avalon_ps2_slave_writedata),   //                   .writedata
		.readdata    (mm_interconnect_0_ps2_port_avalon_ps2_slave_readdata),    //                   .readdata
		.waitrequest (mm_interconnect_0_ps2_port_avalon_ps2_slave_waitrequest), //                   .waitrequest
		.irq         (irq_mapper_receiver1_irq),                                //          interrupt.irq
		.PS2_CLK     (ps2_port_CLK),                                            // external_interface.export
		.PS2_DAT     (ps2_port_DAT)                                             //                   .export
	);

	Computer_System_PS2_Port ps2_port_dual (
		.clk         (system_pll_sys_clk_clk),                                       //                clk.clk
		.reset       (rst_controller_reset_out_reset),                               //              reset.reset
		.address     (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_address),     //   avalon_ps2_slave.address
		.chipselect  (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_chipselect),  //                   .chipselect
		.byteenable  (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_byteenable),  //                   .byteenable
		.read        (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_read),        //                   .read
		.write       (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_write),       //                   .write
		.writedata   (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_writedata),   //                   .writedata
		.readdata    (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_readdata),    //                   .readdata
		.waitrequest (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_waitrequest), //                   .waitrequest
		.irq         (irq_mapper_receiver2_irq),                                     //          interrupt.irq
		.PS2_CLK     (ps2_port_dual_CLK),                                            // external_interface.export
		.PS2_DAT     (ps2_port_dual_DAT)                                             //                   .export
	);

	altera_up_avalon_video_dma_ctrl_addr_trans #(
		.ADDRESS_TRANSLATION_MASK (32'b11000000000000000000000000000000)
	) pixel_dma_addr_translation (
		.clk                (system_pll_sys_clk_clk),                                         //  clock.clk
		.reset              (rst_controller_reset_out_reset),                                 //  reset.reset
		.slave_address      (mm_interconnect_0_pixel_dma_addr_translation_slave_address),     //  slave.address
		.slave_byteenable   (mm_interconnect_0_pixel_dma_addr_translation_slave_byteenable),  //       .byteenable
		.slave_read         (mm_interconnect_0_pixel_dma_addr_translation_slave_read),        //       .read
		.slave_write        (mm_interconnect_0_pixel_dma_addr_translation_slave_write),       //       .write
		.slave_writedata    (mm_interconnect_0_pixel_dma_addr_translation_slave_writedata),   //       .writedata
		.slave_readdata     (mm_interconnect_0_pixel_dma_addr_translation_slave_readdata),    //       .readdata
		.slave_waitrequest  (mm_interconnect_0_pixel_dma_addr_translation_slave_waitrequest), //       .waitrequest
		.master_readdata    (pixel_dma_addr_translation_master_readdata),                     // master.readdata
		.master_waitrequest (pixel_dma_addr_translation_master_waitrequest),                  //       .waitrequest
		.master_address     (pixel_dma_addr_translation_master_address),                      //       .address
		.master_byteenable  (pixel_dma_addr_translation_master_byteenable),                   //       .byteenable
		.master_read        (pixel_dma_addr_translation_master_read),                         //       .read
		.master_write       (pixel_dma_addr_translation_master_write),                        //       .write
		.master_writedata   (pixel_dma_addr_translation_master_writedata)                     //       .writedata
	);

	Computer_System_Pushbuttons pushbuttons (
		.clk        (system_pll_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_pushbuttons_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pushbuttons_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pushbuttons_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pushbuttons_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pushbuttons_s1_readdata),   //                    .readdata
		.in_port    (pushbuttons_export),                          // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                     //                 irq.irq
	);

	Computer_System_SDRAM sdram (
		.clk            (system_pll_sys_clk_clk),                   //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	Computer_System_Slider_Switches slider_switches (
		.clk      (system_pll_sys_clk_clk),                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_slider_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_slider_switches_s1_readdata), //                    .readdata
		.in_port  (slider_switches_export)                         // external_connection.export
	);

	Computer_System_SysID sysid (
		.clock    (system_pll_sys_clk_clk),                         //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	Computer_System_System_PLL system_pll (
		.ref_clk_clk        (system_pll_ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (system_pll_ref_reset_reset),    //    ref_reset.reset
		.sys_clk_clk        (system_pll_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                 //    sdram_clk.clk
		.reset_source_reset (system_pll_reset_source_reset)  // reset_source.reset
	);

	Computer_System_VGA_Subsystem vga_subsystem (
		.char_buffer_control_slave_address    (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_address),    // char_buffer_control_slave.address
		.char_buffer_control_slave_byteenable (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_byteenable), //                          .byteenable
		.char_buffer_control_slave_read       (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_read),       //                          .read
		.char_buffer_control_slave_write      (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_write),      //                          .write
		.char_buffer_control_slave_writedata  (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_writedata),  //                          .writedata
		.char_buffer_control_slave_readdata   (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_readdata),   //                          .readdata
		.char_buffer_slave_address            (mm_interconnect_0_vga_subsystem_char_buffer_slave_address),            //         char_buffer_slave.address
		.char_buffer_slave_clken              (mm_interconnect_0_vga_subsystem_char_buffer_slave_clken),              //                          .clken
		.char_buffer_slave_chipselect         (mm_interconnect_0_vga_subsystem_char_buffer_slave_chipselect),         //                          .chipselect
		.char_buffer_slave_write              (mm_interconnect_0_vga_subsystem_char_buffer_slave_write),              //                          .write
		.char_buffer_slave_readdata           (mm_interconnect_0_vga_subsystem_char_buffer_slave_readdata),           //                          .readdata
		.char_buffer_slave_writedata          (mm_interconnect_0_vga_subsystem_char_buffer_slave_writedata),          //                          .writedata
		.char_buffer_slave_byteenable         (mm_interconnect_0_vga_subsystem_char_buffer_slave_byteenable),         //                          .byteenable
		.pixel_dma_control_slave_address      (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_address),      //   pixel_dma_control_slave.address
		.pixel_dma_control_slave_byteenable   (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_byteenable),   //                          .byteenable
		.pixel_dma_control_slave_read         (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_read),         //                          .read
		.pixel_dma_control_slave_write        (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_write),        //                          .write
		.pixel_dma_control_slave_writedata    (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_writedata),    //                          .writedata
		.pixel_dma_control_slave_readdata     (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_readdata),     //                          .readdata
		.pixel_dma_master_address             (vga_subsystem_pixel_dma_master_address),                               //          pixel_dma_master.address
		.pixel_dma_master_waitrequest         (vga_subsystem_pixel_dma_master_waitrequest),                           //                          .waitrequest
		.pixel_dma_master_lock                (vga_subsystem_pixel_dma_master_lock),                                  //                          .lock
		.pixel_dma_master_read                (vga_subsystem_pixel_dma_master_read),                                  //                          .read
		.pixel_dma_master_readdata            (vga_subsystem_pixel_dma_master_readdata),                              //                          .readdata
		.pixel_dma_master_readdatavalid       (vga_subsystem_pixel_dma_master_readdatavalid),                         //                          .readdatavalid
		.rgb_slave_read                       (mm_interconnect_0_vga_subsystem_rgb_slave_read),                       //                 rgb_slave.read
		.rgb_slave_readdata                   (mm_interconnect_0_vga_subsystem_rgb_slave_readdata),                   //                          .readdata
		.sys_clk_clk                          (system_pll_sys_clk_clk),                                               //                   sys_clk.clk
		.sys_reset_reset_n                    (~rst_controller_006_reset_out_reset),                                  //                 sys_reset.reset_n
		.vga_CLK                              (vga_CLK),                                                              //                       vga.CLK
		.vga_HS                               (vga_HS),                                                               //                          .HS
		.vga_VS                               (vga_VS),                                                               //                          .VS
		.vga_BLANK                            (vga_BLANK),                                                            //                          .BLANK
		.vga_SYNC                             (vga_SYNC),                                                             //                          .SYNC
		.vga_R                                (vga_R),                                                                //                          .R
		.vga_G                                (vga_G),                                                                //                          .G
		.vga_B                                (vga_B),                                                                //                          .B
		.vga_clk_clk                          (video_pll_vga_clk_clk),                                                //                   vga_clk.clk
		.vga_reset_reset_n                    (~video_pll_reset_source_reset)                                         //                 vga_reset.reset_n
	);

	altera_up_avalon_video_dma_ctrl_addr_trans #(
		.ADDRESS_TRANSLATION_MASK (32'b11000000000000000000000000000000)
	) video_in_dma_addr_translation (
		.clk                (system_pll_sys_clk_clk),                                            //  clock.clk
		.reset              (rst_controller_reset_out_reset),                                    //  reset.reset
		.slave_address      (mm_interconnect_0_video_in_dma_addr_translation_slave_address),     //  slave.address
		.slave_byteenable   (mm_interconnect_0_video_in_dma_addr_translation_slave_byteenable),  //       .byteenable
		.slave_read         (mm_interconnect_0_video_in_dma_addr_translation_slave_read),        //       .read
		.slave_write        (mm_interconnect_0_video_in_dma_addr_translation_slave_write),       //       .write
		.slave_writedata    (mm_interconnect_0_video_in_dma_addr_translation_slave_writedata),   //       .writedata
		.slave_readdata     (mm_interconnect_0_video_in_dma_addr_translation_slave_readdata),    //       .readdata
		.slave_waitrequest  (mm_interconnect_0_video_in_dma_addr_translation_slave_waitrequest), //       .waitrequest
		.master_readdata    (video_in_dma_addr_translation_master_readdata),                     // master.readdata
		.master_waitrequest (video_in_dma_addr_translation_master_waitrequest),                  //       .waitrequest
		.master_address     (video_in_dma_addr_translation_master_address),                      //       .address
		.master_byteenable  (video_in_dma_addr_translation_master_byteenable),                   //       .byteenable
		.master_read        (video_in_dma_addr_translation_master_read),                         //       .read
		.master_write       (video_in_dma_addr_translation_master_write),                        //       .write
		.master_writedata   (video_in_dma_addr_translation_master_writedata)                     //       .writedata
	);

	Computer_System_Video_In_Subsystem video_in_subsystem (
		.sys_clk_clk                                      (system_pll_sys_clk_clk),                                                                //                               sys_clk.clk
		.sys_reset_reset_n                                (~rst_controller_007_reset_out_reset),                                                   //                             sys_reset.reset_n
		.video_in_TD_CLK27                                (video_in_TD_CLK27),                                                                     //                              video_in.TD_CLK27
		.video_in_TD_DATA                                 (video_in_TD_DATA),                                                                      //                                      .TD_DATA
		.video_in_TD_HS                                   (video_in_TD_HS),                                                                        //                                      .TD_HS
		.video_in_TD_VS                                   (video_in_TD_VS),                                                                        //                                      .TD_VS
		.video_in_clk27_reset                             (video_in_clk27_reset),                                                                  //                                      .clk27_reset
		.video_in_TD_RESET                                (video_in_TD_RESET),                                                                     //                                      .TD_RESET
		.video_in_overflow_flag                           (video_in_overflow_flag),                                                                //                                      .overflow_flag
		.video_in_dma_control_slave_address               (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_address),               //            video_in_dma_control_slave.address
		.video_in_dma_control_slave_byteenable            (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_byteenable),            //                                      .byteenable
		.video_in_dma_control_slave_read                  (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_read),                  //                                      .read
		.video_in_dma_control_slave_write                 (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_write),                 //                                      .write
		.video_in_dma_control_slave_writedata             (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_writedata),             //                                      .writedata
		.video_in_dma_control_slave_readdata              (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_readdata),              //                                      .readdata
		.video_in_dma_master_address                      (video_in_subsystem_video_in_dma_master_address),                                        //                   video_in_dma_master.address
		.video_in_dma_master_waitrequest                  (video_in_subsystem_video_in_dma_master_waitrequest),                                    //                                      .waitrequest
		.video_in_dma_master_write                        (video_in_subsystem_video_in_dma_master_write),                                          //                                      .write
		.video_in_dma_master_writedata                    (video_in_subsystem_video_in_dma_master_writedata),                                      //                                      .writedata
		.video_in_edge_detection_control_slave_address    (mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_address),    // video_in_edge_detection_control_slave.address
		.video_in_edge_detection_control_slave_write_n    (~mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_write),     //                                      .write_n
		.video_in_edge_detection_control_slave_writedata  (mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_writedata),  //                                      .writedata
		.video_in_edge_detection_control_slave_chipselect (mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_chipselect), //                                      .chipselect
		.video_in_edge_detection_control_slave_readdata   (mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_readdata)    //                                      .readdata
	);

	Computer_System_Video_PLL video_pll (
		.ref_clk_clk        (video_pll_ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (video_pll_ref_reset_reset),    //    ref_reset.reset
		.vga_clk_clk        (video_pll_vga_clk_clk),        //      vga_clk.clk
		.reset_source_reset (video_pll_reset_source_reset)  // reset_source.reset
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) nios2_custom_instruction_master_translator (
		.ci_slave_result           (),                                                                     //        ci_slave.result
		.ci_slave_multi_clk        (nios2_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios2_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios2_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios2_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios2_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios2_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (nios2_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (nios2_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (nios2_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (nios2_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (nios2_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (nios2_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (nios2_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (nios2_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (nios2_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (nios2_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_result     (),                                                                     //  comb_ci_master.result
		.multi_ci_master_clk       (nios2_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios2_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios2_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios2_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios2_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios2_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios2_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios2_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios2_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios2_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios2_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios2_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios2_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios2_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios2_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios2_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_dataa            (32'b00000000000000000000000000000000),                                 //     (terminated)
		.ci_slave_datab            (32'b00000000000000000000000000000000),                                 //     (terminated)
		.ci_slave_n                (8'b00000000),                                                          //     (terminated)
		.ci_slave_readra           (1'b0),                                                                 //     (terminated)
		.ci_slave_readrb           (1'b0),                                                                 //     (terminated)
		.ci_slave_writerc          (1'b0),                                                                 //     (terminated)
		.ci_slave_a                (5'b00000),                                                             //     (terminated)
		.ci_slave_b                (5'b00000),                                                             //     (terminated)
		.ci_slave_c                (5'b00000),                                                             //     (terminated)
		.ci_slave_ipending         (32'b00000000000000000000000000000000),                                 //     (terminated)
		.ci_slave_estatus          (1'b0),                                                                 //     (terminated)
		.comb_ci_master_dataa      (),                                                                     //     (terminated)
		.comb_ci_master_datab      (),                                                                     //     (terminated)
		.comb_ci_master_n          (),                                                                     //     (terminated)
		.comb_ci_master_readra     (),                                                                     //     (terminated)
		.comb_ci_master_readrb     (),                                                                     //     (terminated)
		.comb_ci_master_writerc    (),                                                                     //     (terminated)
		.comb_ci_master_a          (),                                                                     //     (terminated)
		.comb_ci_master_b          (),                                                                     //     (terminated)
		.comb_ci_master_c          (),                                                                     //     (terminated)
		.comb_ci_master_ipending   (),                                                                     //     (terminated)
		.comb_ci_master_estatus    ()                                                                      //     (terminated)
	);

	Computer_System_Nios2_custom_instruction_master_multi_xconnect nios2_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios2_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios2_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios2_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios2_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios2_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios2_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios2_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios2_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios2_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios2_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                     //           .ipending
		.ci_slave_estatus     (),                                                                     //           .estatus
		.ci_slave_clk         (nios2_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios2_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios2_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios2_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios2_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios2_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios2_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios2_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios2_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios2_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios2_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios2_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios2_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios2_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios2_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios2_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios2_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios2_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios2_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios2_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (2),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) nios2_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios2_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (nios2_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (nios2_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (nios2_custom_instruction_master_multi_slave_translator0_ci_master_n),      //          .n
		.ci_master_clk       (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (nios2_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_readra    (),                                                                         // (terminated)
		.ci_master_readrb    (),                                                                         // (terminated)
		.ci_master_writerc   (),                                                                         // (terminated)
		.ci_master_a         (),                                                                         // (terminated)
		.ci_master_b         (),                                                                         // (terminated)
		.ci_master_c         (),                                                                         // (terminated)
		.ci_master_ipending  (),                                                                         // (terminated)
		.ci_master_estatus   (),                                                                         // (terminated)
		.ci_master_reset_req ()                                                                          // (terminated)
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) nios2_2nd_core_custom_instruction_master_translator (
		.ci_slave_result           (),                                                                              //        ci_slave.result
		.ci_slave_multi_clk        (nios2_2nd_core_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios2_2nd_core_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios2_2nd_core_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios2_2nd_core_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios2_2nd_core_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios2_2nd_core_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (nios2_2nd_core_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (nios2_2nd_core_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (nios2_2nd_core_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (nios2_2nd_core_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (nios2_2nd_core_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (nios2_2nd_core_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (nios2_2nd_core_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (nios2_2nd_core_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (nios2_2nd_core_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (nios2_2nd_core_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_result     (),                                                                              //  comb_ci_master.result
		.multi_ci_master_clk       (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_dataa            (32'b00000000000000000000000000000000),                                          //     (terminated)
		.ci_slave_datab            (32'b00000000000000000000000000000000),                                          //     (terminated)
		.ci_slave_n                (8'b00000000),                                                                   //     (terminated)
		.ci_slave_readra           (1'b0),                                                                          //     (terminated)
		.ci_slave_readrb           (1'b0),                                                                          //     (terminated)
		.ci_slave_writerc          (1'b0),                                                                          //     (terminated)
		.ci_slave_a                (5'b00000),                                                                      //     (terminated)
		.ci_slave_b                (5'b00000),                                                                      //     (terminated)
		.ci_slave_c                (5'b00000),                                                                      //     (terminated)
		.ci_slave_ipending         (32'b00000000000000000000000000000000),                                          //     (terminated)
		.ci_slave_estatus          (1'b0),                                                                          //     (terminated)
		.comb_ci_master_dataa      (),                                                                              //     (terminated)
		.comb_ci_master_datab      (),                                                                              //     (terminated)
		.comb_ci_master_n          (),                                                                              //     (terminated)
		.comb_ci_master_readra     (),                                                                              //     (terminated)
		.comb_ci_master_readrb     (),                                                                              //     (terminated)
		.comb_ci_master_writerc    (),                                                                              //     (terminated)
		.comb_ci_master_a          (),                                                                              //     (terminated)
		.comb_ci_master_b          (),                                                                              //     (terminated)
		.comb_ci_master_c          (),                                                                              //     (terminated)
		.comb_ci_master_ipending   (),                                                                              //     (terminated)
		.comb_ci_master_estatus    ()                                                                               //     (terminated)
	);

	Computer_System_Nios2_custom_instruction_master_multi_xconnect nios2_2nd_core_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                              //           .ipending
		.ci_slave_estatus     (),                                                                              //           .estatus
		.ci_slave_clk         (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (2),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) nios2_2nd_core_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_n),      //          .n
		.ci_master_clk       (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_readra    (),                                                                                  // (terminated)
		.ci_master_readrb    (),                                                                                  // (terminated)
		.ci_master_writerc   (),                                                                                  // (terminated)
		.ci_master_a         (),                                                                                  // (terminated)
		.ci_master_b         (),                                                                                  // (terminated)
		.ci_master_c         (),                                                                                  // (terminated)
		.ci_master_ipending  (),                                                                                  // (terminated)
		.ci_master_estatus   (),                                                                                  // (terminated)
		.ci_master_reset_req ()                                                                                   // (terminated)
	);

	Computer_System_mm_interconnect_0 mm_interconnect_0 (
		.ARM_A9_HPS_h2f_axi_master_awid                                           (arm_a9_hps_h2f_axi_master_awid),                                                        //                                          ARM_A9_HPS_h2f_axi_master.awid
		.ARM_A9_HPS_h2f_axi_master_awaddr                                         (arm_a9_hps_h2f_axi_master_awaddr),                                                      //                                                                   .awaddr
		.ARM_A9_HPS_h2f_axi_master_awlen                                          (arm_a9_hps_h2f_axi_master_awlen),                                                       //                                                                   .awlen
		.ARM_A9_HPS_h2f_axi_master_awsize                                         (arm_a9_hps_h2f_axi_master_awsize),                                                      //                                                                   .awsize
		.ARM_A9_HPS_h2f_axi_master_awburst                                        (arm_a9_hps_h2f_axi_master_awburst),                                                     //                                                                   .awburst
		.ARM_A9_HPS_h2f_axi_master_awlock                                         (arm_a9_hps_h2f_axi_master_awlock),                                                      //                                                                   .awlock
		.ARM_A9_HPS_h2f_axi_master_awcache                                        (arm_a9_hps_h2f_axi_master_awcache),                                                     //                                                                   .awcache
		.ARM_A9_HPS_h2f_axi_master_awprot                                         (arm_a9_hps_h2f_axi_master_awprot),                                                      //                                                                   .awprot
		.ARM_A9_HPS_h2f_axi_master_awvalid                                        (arm_a9_hps_h2f_axi_master_awvalid),                                                     //                                                                   .awvalid
		.ARM_A9_HPS_h2f_axi_master_awready                                        (arm_a9_hps_h2f_axi_master_awready),                                                     //                                                                   .awready
		.ARM_A9_HPS_h2f_axi_master_wid                                            (arm_a9_hps_h2f_axi_master_wid),                                                         //                                                                   .wid
		.ARM_A9_HPS_h2f_axi_master_wdata                                          (arm_a9_hps_h2f_axi_master_wdata),                                                       //                                                                   .wdata
		.ARM_A9_HPS_h2f_axi_master_wstrb                                          (arm_a9_hps_h2f_axi_master_wstrb),                                                       //                                                                   .wstrb
		.ARM_A9_HPS_h2f_axi_master_wlast                                          (arm_a9_hps_h2f_axi_master_wlast),                                                       //                                                                   .wlast
		.ARM_A9_HPS_h2f_axi_master_wvalid                                         (arm_a9_hps_h2f_axi_master_wvalid),                                                      //                                                                   .wvalid
		.ARM_A9_HPS_h2f_axi_master_wready                                         (arm_a9_hps_h2f_axi_master_wready),                                                      //                                                                   .wready
		.ARM_A9_HPS_h2f_axi_master_bid                                            (arm_a9_hps_h2f_axi_master_bid),                                                         //                                                                   .bid
		.ARM_A9_HPS_h2f_axi_master_bresp                                          (arm_a9_hps_h2f_axi_master_bresp),                                                       //                                                                   .bresp
		.ARM_A9_HPS_h2f_axi_master_bvalid                                         (arm_a9_hps_h2f_axi_master_bvalid),                                                      //                                                                   .bvalid
		.ARM_A9_HPS_h2f_axi_master_bready                                         (arm_a9_hps_h2f_axi_master_bready),                                                      //                                                                   .bready
		.ARM_A9_HPS_h2f_axi_master_arid                                           (arm_a9_hps_h2f_axi_master_arid),                                                        //                                                                   .arid
		.ARM_A9_HPS_h2f_axi_master_araddr                                         (arm_a9_hps_h2f_axi_master_araddr),                                                      //                                                                   .araddr
		.ARM_A9_HPS_h2f_axi_master_arlen                                          (arm_a9_hps_h2f_axi_master_arlen),                                                       //                                                                   .arlen
		.ARM_A9_HPS_h2f_axi_master_arsize                                         (arm_a9_hps_h2f_axi_master_arsize),                                                      //                                                                   .arsize
		.ARM_A9_HPS_h2f_axi_master_arburst                                        (arm_a9_hps_h2f_axi_master_arburst),                                                     //                                                                   .arburst
		.ARM_A9_HPS_h2f_axi_master_arlock                                         (arm_a9_hps_h2f_axi_master_arlock),                                                      //                                                                   .arlock
		.ARM_A9_HPS_h2f_axi_master_arcache                                        (arm_a9_hps_h2f_axi_master_arcache),                                                     //                                                                   .arcache
		.ARM_A9_HPS_h2f_axi_master_arprot                                         (arm_a9_hps_h2f_axi_master_arprot),                                                      //                                                                   .arprot
		.ARM_A9_HPS_h2f_axi_master_arvalid                                        (arm_a9_hps_h2f_axi_master_arvalid),                                                     //                                                                   .arvalid
		.ARM_A9_HPS_h2f_axi_master_arready                                        (arm_a9_hps_h2f_axi_master_arready),                                                     //                                                                   .arready
		.ARM_A9_HPS_h2f_axi_master_rid                                            (arm_a9_hps_h2f_axi_master_rid),                                                         //                                                                   .rid
		.ARM_A9_HPS_h2f_axi_master_rdata                                          (arm_a9_hps_h2f_axi_master_rdata),                                                       //                                                                   .rdata
		.ARM_A9_HPS_h2f_axi_master_rresp                                          (arm_a9_hps_h2f_axi_master_rresp),                                                       //                                                                   .rresp
		.ARM_A9_HPS_h2f_axi_master_rlast                                          (arm_a9_hps_h2f_axi_master_rlast),                                                       //                                                                   .rlast
		.ARM_A9_HPS_h2f_axi_master_rvalid                                         (arm_a9_hps_h2f_axi_master_rvalid),                                                      //                                                                   .rvalid
		.ARM_A9_HPS_h2f_axi_master_rready                                         (arm_a9_hps_h2f_axi_master_rready),                                                      //                                                                   .rready
		.ARM_A9_HPS_h2f_lw_axi_master_awid                                        (arm_a9_hps_h2f_lw_axi_master_awid),                                                     //                                       ARM_A9_HPS_h2f_lw_axi_master.awid
		.ARM_A9_HPS_h2f_lw_axi_master_awaddr                                      (arm_a9_hps_h2f_lw_axi_master_awaddr),                                                   //                                                                   .awaddr
		.ARM_A9_HPS_h2f_lw_axi_master_awlen                                       (arm_a9_hps_h2f_lw_axi_master_awlen),                                                    //                                                                   .awlen
		.ARM_A9_HPS_h2f_lw_axi_master_awsize                                      (arm_a9_hps_h2f_lw_axi_master_awsize),                                                   //                                                                   .awsize
		.ARM_A9_HPS_h2f_lw_axi_master_awburst                                     (arm_a9_hps_h2f_lw_axi_master_awburst),                                                  //                                                                   .awburst
		.ARM_A9_HPS_h2f_lw_axi_master_awlock                                      (arm_a9_hps_h2f_lw_axi_master_awlock),                                                   //                                                                   .awlock
		.ARM_A9_HPS_h2f_lw_axi_master_awcache                                     (arm_a9_hps_h2f_lw_axi_master_awcache),                                                  //                                                                   .awcache
		.ARM_A9_HPS_h2f_lw_axi_master_awprot                                      (arm_a9_hps_h2f_lw_axi_master_awprot),                                                   //                                                                   .awprot
		.ARM_A9_HPS_h2f_lw_axi_master_awvalid                                     (arm_a9_hps_h2f_lw_axi_master_awvalid),                                                  //                                                                   .awvalid
		.ARM_A9_HPS_h2f_lw_axi_master_awready                                     (arm_a9_hps_h2f_lw_axi_master_awready),                                                  //                                                                   .awready
		.ARM_A9_HPS_h2f_lw_axi_master_wid                                         (arm_a9_hps_h2f_lw_axi_master_wid),                                                      //                                                                   .wid
		.ARM_A9_HPS_h2f_lw_axi_master_wdata                                       (arm_a9_hps_h2f_lw_axi_master_wdata),                                                    //                                                                   .wdata
		.ARM_A9_HPS_h2f_lw_axi_master_wstrb                                       (arm_a9_hps_h2f_lw_axi_master_wstrb),                                                    //                                                                   .wstrb
		.ARM_A9_HPS_h2f_lw_axi_master_wlast                                       (arm_a9_hps_h2f_lw_axi_master_wlast),                                                    //                                                                   .wlast
		.ARM_A9_HPS_h2f_lw_axi_master_wvalid                                      (arm_a9_hps_h2f_lw_axi_master_wvalid),                                                   //                                                                   .wvalid
		.ARM_A9_HPS_h2f_lw_axi_master_wready                                      (arm_a9_hps_h2f_lw_axi_master_wready),                                                   //                                                                   .wready
		.ARM_A9_HPS_h2f_lw_axi_master_bid                                         (arm_a9_hps_h2f_lw_axi_master_bid),                                                      //                                                                   .bid
		.ARM_A9_HPS_h2f_lw_axi_master_bresp                                       (arm_a9_hps_h2f_lw_axi_master_bresp),                                                    //                                                                   .bresp
		.ARM_A9_HPS_h2f_lw_axi_master_bvalid                                      (arm_a9_hps_h2f_lw_axi_master_bvalid),                                                   //                                                                   .bvalid
		.ARM_A9_HPS_h2f_lw_axi_master_bready                                      (arm_a9_hps_h2f_lw_axi_master_bready),                                                   //                                                                   .bready
		.ARM_A9_HPS_h2f_lw_axi_master_arid                                        (arm_a9_hps_h2f_lw_axi_master_arid),                                                     //                                                                   .arid
		.ARM_A9_HPS_h2f_lw_axi_master_araddr                                      (arm_a9_hps_h2f_lw_axi_master_araddr),                                                   //                                                                   .araddr
		.ARM_A9_HPS_h2f_lw_axi_master_arlen                                       (arm_a9_hps_h2f_lw_axi_master_arlen),                                                    //                                                                   .arlen
		.ARM_A9_HPS_h2f_lw_axi_master_arsize                                      (arm_a9_hps_h2f_lw_axi_master_arsize),                                                   //                                                                   .arsize
		.ARM_A9_HPS_h2f_lw_axi_master_arburst                                     (arm_a9_hps_h2f_lw_axi_master_arburst),                                                  //                                                                   .arburst
		.ARM_A9_HPS_h2f_lw_axi_master_arlock                                      (arm_a9_hps_h2f_lw_axi_master_arlock),                                                   //                                                                   .arlock
		.ARM_A9_HPS_h2f_lw_axi_master_arcache                                     (arm_a9_hps_h2f_lw_axi_master_arcache),                                                  //                                                                   .arcache
		.ARM_A9_HPS_h2f_lw_axi_master_arprot                                      (arm_a9_hps_h2f_lw_axi_master_arprot),                                                   //                                                                   .arprot
		.ARM_A9_HPS_h2f_lw_axi_master_arvalid                                     (arm_a9_hps_h2f_lw_axi_master_arvalid),                                                  //                                                                   .arvalid
		.ARM_A9_HPS_h2f_lw_axi_master_arready                                     (arm_a9_hps_h2f_lw_axi_master_arready),                                                  //                                                                   .arready
		.ARM_A9_HPS_h2f_lw_axi_master_rid                                         (arm_a9_hps_h2f_lw_axi_master_rid),                                                      //                                                                   .rid
		.ARM_A9_HPS_h2f_lw_axi_master_rdata                                       (arm_a9_hps_h2f_lw_axi_master_rdata),                                                    //                                                                   .rdata
		.ARM_A9_HPS_h2f_lw_axi_master_rresp                                       (arm_a9_hps_h2f_lw_axi_master_rresp),                                                    //                                                                   .rresp
		.ARM_A9_HPS_h2f_lw_axi_master_rlast                                       (arm_a9_hps_h2f_lw_axi_master_rlast),                                                    //                                                                   .rlast
		.ARM_A9_HPS_h2f_lw_axi_master_rvalid                                      (arm_a9_hps_h2f_lw_axi_master_rvalid),                                                   //                                                                   .rvalid
		.ARM_A9_HPS_h2f_lw_axi_master_rready                                      (arm_a9_hps_h2f_lw_axi_master_rready),                                                   //                                                                   .rready
		.System_PLL_sys_clk_clk                                                   (system_pll_sys_clk_clk),                                                                //                                                 System_PLL_sys_clk.clk
		.ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_008_reset_out_reset),                                                    // ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset                (rst_controller_reset_out_reset),                                                        //                JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset.reset
		.Nios2_2nd_Core_reset_reset_bridge_in_reset_reset                         (rst_controller_005_reset_out_reset),                                                    //                         Nios2_2nd_Core_reset_reset_bridge_in_reset.reset
		.Nios2_reset_reset_bridge_in_reset_reset                                  (rst_controller_004_reset_out_reset),                                                    //                                  Nios2_reset_reset_bridge_in_reset.reset
		.Video_In_DMA_Addr_Translation_reset_reset_bridge_in_reset_reset          (rst_controller_reset_out_reset),                                                        //          Video_In_DMA_Addr_Translation_reset_reset_bridge_in_reset.reset
		.Char_DMA_Addr_Translation_master_address                                 (char_dma_addr_translation_master_address),                                              //                                   Char_DMA_Addr_Translation_master.address
		.Char_DMA_Addr_Translation_master_waitrequest                             (char_dma_addr_translation_master_waitrequest),                                          //                                                                   .waitrequest
		.Char_DMA_Addr_Translation_master_byteenable                              (char_dma_addr_translation_master_byteenable),                                           //                                                                   .byteenable
		.Char_DMA_Addr_Translation_master_read                                    (char_dma_addr_translation_master_read),                                                 //                                                                   .read
		.Char_DMA_Addr_Translation_master_readdata                                (char_dma_addr_translation_master_readdata),                                             //                                                                   .readdata
		.Char_DMA_Addr_Translation_master_write                                   (char_dma_addr_translation_master_write),                                                //                                                                   .write
		.Char_DMA_Addr_Translation_master_writedata                               (char_dma_addr_translation_master_writedata),                                            //                                                                   .writedata
		.JTAG_to_FPGA_Bridge_master_address                                       (jtag_to_fpga_bridge_master_address),                                                    //                                         JTAG_to_FPGA_Bridge_master.address
		.JTAG_to_FPGA_Bridge_master_waitrequest                                   (jtag_to_fpga_bridge_master_waitrequest),                                                //                                                                   .waitrequest
		.JTAG_to_FPGA_Bridge_master_byteenable                                    (jtag_to_fpga_bridge_master_byteenable),                                                 //                                                                   .byteenable
		.JTAG_to_FPGA_Bridge_master_read                                          (jtag_to_fpga_bridge_master_read),                                                       //                                                                   .read
		.JTAG_to_FPGA_Bridge_master_readdata                                      (jtag_to_fpga_bridge_master_readdata),                                                   //                                                                   .readdata
		.JTAG_to_FPGA_Bridge_master_readdatavalid                                 (jtag_to_fpga_bridge_master_readdatavalid),                                              //                                                                   .readdatavalid
		.JTAG_to_FPGA_Bridge_master_write                                         (jtag_to_fpga_bridge_master_write),                                                      //                                                                   .write
		.JTAG_to_FPGA_Bridge_master_writedata                                     (jtag_to_fpga_bridge_master_writedata),                                                  //                                                                   .writedata
		.Nios2_data_master_address                                                (nios2_data_master_address),                                                             //                                                  Nios2_data_master.address
		.Nios2_data_master_waitrequest                                            (nios2_data_master_waitrequest),                                                         //                                                                   .waitrequest
		.Nios2_data_master_byteenable                                             (nios2_data_master_byteenable),                                                          //                                                                   .byteenable
		.Nios2_data_master_read                                                   (nios2_data_master_read),                                                                //                                                                   .read
		.Nios2_data_master_readdata                                               (nios2_data_master_readdata),                                                            //                                                                   .readdata
		.Nios2_data_master_write                                                  (nios2_data_master_write),                                                               //                                                                   .write
		.Nios2_data_master_writedata                                              (nios2_data_master_writedata),                                                           //                                                                   .writedata
		.Nios2_data_master_debugaccess                                            (nios2_data_master_debugaccess),                                                         //                                                                   .debugaccess
		.Nios2_instruction_master_address                                         (nios2_instruction_master_address),                                                      //                                           Nios2_instruction_master.address
		.Nios2_instruction_master_waitrequest                                     (nios2_instruction_master_waitrequest),                                                  //                                                                   .waitrequest
		.Nios2_instruction_master_read                                            (nios2_instruction_master_read),                                                         //                                                                   .read
		.Nios2_instruction_master_readdata                                        (nios2_instruction_master_readdata),                                                     //                                                                   .readdata
		.Nios2_instruction_master_readdatavalid                                   (nios2_instruction_master_readdatavalid),                                                //                                                                   .readdatavalid
		.Nios2_2nd_Core_data_master_address                                       (nios2_2nd_core_data_master_address),                                                    //                                         Nios2_2nd_Core_data_master.address
		.Nios2_2nd_Core_data_master_waitrequest                                   (nios2_2nd_core_data_master_waitrequest),                                                //                                                                   .waitrequest
		.Nios2_2nd_Core_data_master_byteenable                                    (nios2_2nd_core_data_master_byteenable),                                                 //                                                                   .byteenable
		.Nios2_2nd_Core_data_master_read                                          (nios2_2nd_core_data_master_read),                                                       //                                                                   .read
		.Nios2_2nd_Core_data_master_readdata                                      (nios2_2nd_core_data_master_readdata),                                                   //                                                                   .readdata
		.Nios2_2nd_Core_data_master_write                                         (nios2_2nd_core_data_master_write),                                                      //                                                                   .write
		.Nios2_2nd_Core_data_master_writedata                                     (nios2_2nd_core_data_master_writedata),                                                  //                                                                   .writedata
		.Nios2_2nd_Core_data_master_debugaccess                                   (nios2_2nd_core_data_master_debugaccess),                                                //                                                                   .debugaccess
		.Nios2_2nd_Core_instruction_master_address                                (nios2_2nd_core_instruction_master_address),                                             //                                  Nios2_2nd_Core_instruction_master.address
		.Nios2_2nd_Core_instruction_master_waitrequest                            (nios2_2nd_core_instruction_master_waitrequest),                                         //                                                                   .waitrequest
		.Nios2_2nd_Core_instruction_master_read                                   (nios2_2nd_core_instruction_master_read),                                                //                                                                   .read
		.Nios2_2nd_Core_instruction_master_readdata                               (nios2_2nd_core_instruction_master_readdata),                                            //                                                                   .readdata
		.Nios2_2nd_Core_instruction_master_readdatavalid                          (nios2_2nd_core_instruction_master_readdatavalid),                                       //                                                                   .readdatavalid
		.Pixel_DMA_Addr_Translation_master_address                                (pixel_dma_addr_translation_master_address),                                             //                                  Pixel_DMA_Addr_Translation_master.address
		.Pixel_DMA_Addr_Translation_master_waitrequest                            (pixel_dma_addr_translation_master_waitrequest),                                         //                                                                   .waitrequest
		.Pixel_DMA_Addr_Translation_master_byteenable                             (pixel_dma_addr_translation_master_byteenable),                                          //                                                                   .byteenable
		.Pixel_DMA_Addr_Translation_master_read                                   (pixel_dma_addr_translation_master_read),                                                //                                                                   .read
		.Pixel_DMA_Addr_Translation_master_readdata                               (pixel_dma_addr_translation_master_readdata),                                            //                                                                   .readdata
		.Pixel_DMA_Addr_Translation_master_write                                  (pixel_dma_addr_translation_master_write),                                               //                                                                   .write
		.Pixel_DMA_Addr_Translation_master_writedata                              (pixel_dma_addr_translation_master_writedata),                                           //                                                                   .writedata
		.VGA_Subsystem_pixel_dma_master_address                                   (vga_subsystem_pixel_dma_master_address),                                                //                                     VGA_Subsystem_pixel_dma_master.address
		.VGA_Subsystem_pixel_dma_master_waitrequest                               (vga_subsystem_pixel_dma_master_waitrequest),                                            //                                                                   .waitrequest
		.VGA_Subsystem_pixel_dma_master_read                                      (vga_subsystem_pixel_dma_master_read),                                                   //                                                                   .read
		.VGA_Subsystem_pixel_dma_master_readdata                                  (vga_subsystem_pixel_dma_master_readdata),                                               //                                                                   .readdata
		.VGA_Subsystem_pixel_dma_master_readdatavalid                             (vga_subsystem_pixel_dma_master_readdatavalid),                                          //                                                                   .readdatavalid
		.VGA_Subsystem_pixel_dma_master_lock                                      (vga_subsystem_pixel_dma_master_lock),                                                   //                                                                   .lock
		.Video_In_DMA_Addr_Translation_master_address                             (video_in_dma_addr_translation_master_address),                                          //                               Video_In_DMA_Addr_Translation_master.address
		.Video_In_DMA_Addr_Translation_master_waitrequest                         (video_in_dma_addr_translation_master_waitrequest),                                      //                                                                   .waitrequest
		.Video_In_DMA_Addr_Translation_master_byteenable                          (video_in_dma_addr_translation_master_byteenable),                                       //                                                                   .byteenable
		.Video_In_DMA_Addr_Translation_master_read                                (video_in_dma_addr_translation_master_read),                                             //                                                                   .read
		.Video_In_DMA_Addr_Translation_master_readdata                            (video_in_dma_addr_translation_master_readdata),                                         //                                                                   .readdata
		.Video_In_DMA_Addr_Translation_master_write                               (video_in_dma_addr_translation_master_write),                                            //                                                                   .write
		.Video_In_DMA_Addr_Translation_master_writedata                           (video_in_dma_addr_translation_master_writedata),                                        //                                                                   .writedata
		.Video_In_Subsystem_video_in_dma_master_address                           (video_in_subsystem_video_in_dma_master_address),                                        //                             Video_In_Subsystem_video_in_dma_master.address
		.Video_In_Subsystem_video_in_dma_master_waitrequest                       (video_in_subsystem_video_in_dma_master_waitrequest),                                    //                                                                   .waitrequest
		.Video_In_Subsystem_video_in_dma_master_write                             (video_in_subsystem_video_in_dma_master_write),                                          //                                                                   .write
		.Video_In_Subsystem_video_in_dma_master_writedata                         (video_in_subsystem_video_in_dma_master_writedata),                                      //                                                                   .writedata
		.ADC_adc_slave_address                                                    (mm_interconnect_0_adc_adc_slave_address),                                               //                                                      ADC_adc_slave.address
		.ADC_adc_slave_write                                                      (mm_interconnect_0_adc_adc_slave_write),                                                 //                                                                   .write
		.ADC_adc_slave_read                                                       (mm_interconnect_0_adc_adc_slave_read),                                                  //                                                                   .read
		.ADC_adc_slave_readdata                                                   (mm_interconnect_0_adc_adc_slave_readdata),                                              //                                                                   .readdata
		.ADC_adc_slave_writedata                                                  (mm_interconnect_0_adc_adc_slave_writedata),                                             //                                                                   .writedata
		.ADC_adc_slave_waitrequest                                                (mm_interconnect_0_adc_adc_slave_waitrequest),                                           //                                                                   .waitrequest
		.Audio_Subsystem_audio_slave_address                                      (mm_interconnect_0_audio_subsystem_audio_slave_address),                                 //                                        Audio_Subsystem_audio_slave.address
		.Audio_Subsystem_audio_slave_write                                        (mm_interconnect_0_audio_subsystem_audio_slave_write),                                   //                                                                   .write
		.Audio_Subsystem_audio_slave_read                                         (mm_interconnect_0_audio_subsystem_audio_slave_read),                                    //                                                                   .read
		.Audio_Subsystem_audio_slave_readdata                                     (mm_interconnect_0_audio_subsystem_audio_slave_readdata),                                //                                                                   .readdata
		.Audio_Subsystem_audio_slave_writedata                                    (mm_interconnect_0_audio_subsystem_audio_slave_writedata),                               //                                                                   .writedata
		.Audio_Subsystem_audio_slave_chipselect                                   (mm_interconnect_0_audio_subsystem_audio_slave_chipselect),                              //                                                                   .chipselect
		.AV_Config_avalon_av_config_slave_address                                 (mm_interconnect_0_av_config_avalon_av_config_slave_address),                            //                                   AV_Config_avalon_av_config_slave.address
		.AV_Config_avalon_av_config_slave_write                                   (mm_interconnect_0_av_config_avalon_av_config_slave_write),                              //                                                                   .write
		.AV_Config_avalon_av_config_slave_read                                    (mm_interconnect_0_av_config_avalon_av_config_slave_read),                               //                                                                   .read
		.AV_Config_avalon_av_config_slave_readdata                                (mm_interconnect_0_av_config_avalon_av_config_slave_readdata),                           //                                                                   .readdata
		.AV_Config_avalon_av_config_slave_writedata                               (mm_interconnect_0_av_config_avalon_av_config_slave_writedata),                          //                                                                   .writedata
		.AV_Config_avalon_av_config_slave_byteenable                              (mm_interconnect_0_av_config_avalon_av_config_slave_byteenable),                         //                                                                   .byteenable
		.AV_Config_avalon_av_config_slave_waitrequest                             (mm_interconnect_0_av_config_avalon_av_config_slave_waitrequest),                        //                                                                   .waitrequest
		.Char_DMA_Addr_Translation_slave_address                                  (mm_interconnect_0_char_dma_addr_translation_slave_address),                             //                                    Char_DMA_Addr_Translation_slave.address
		.Char_DMA_Addr_Translation_slave_write                                    (mm_interconnect_0_char_dma_addr_translation_slave_write),                               //                                                                   .write
		.Char_DMA_Addr_Translation_slave_read                                     (mm_interconnect_0_char_dma_addr_translation_slave_read),                                //                                                                   .read
		.Char_DMA_Addr_Translation_slave_readdata                                 (mm_interconnect_0_char_dma_addr_translation_slave_readdata),                            //                                                                   .readdata
		.Char_DMA_Addr_Translation_slave_writedata                                (mm_interconnect_0_char_dma_addr_translation_slave_writedata),                           //                                                                   .writedata
		.Char_DMA_Addr_Translation_slave_byteenable                               (mm_interconnect_0_char_dma_addr_translation_slave_byteenable),                          //                                                                   .byteenable
		.Char_DMA_Addr_Translation_slave_waitrequest                              (mm_interconnect_0_char_dma_addr_translation_slave_waitrequest),                         //                                                                   .waitrequest
		.Expansion_JP1_s1_address                                                 (mm_interconnect_0_expansion_jp1_s1_address),                                            //                                                   Expansion_JP1_s1.address
		.Expansion_JP1_s1_write                                                   (mm_interconnect_0_expansion_jp1_s1_write),                                              //                                                                   .write
		.Expansion_JP1_s1_readdata                                                (mm_interconnect_0_expansion_jp1_s1_readdata),                                           //                                                                   .readdata
		.Expansion_JP1_s1_writedata                                               (mm_interconnect_0_expansion_jp1_s1_writedata),                                          //                                                                   .writedata
		.Expansion_JP1_s1_chipselect                                              (mm_interconnect_0_expansion_jp1_s1_chipselect),                                         //                                                                   .chipselect
		.F2H_Mem_Window_00000000_windowed_slave_address                           (mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_address),                      //                             F2H_Mem_Window_00000000_windowed_slave.address
		.F2H_Mem_Window_00000000_windowed_slave_write                             (mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_write),                        //                                                                   .write
		.F2H_Mem_Window_00000000_windowed_slave_read                              (mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_read),                         //                                                                   .read
		.F2H_Mem_Window_00000000_windowed_slave_readdata                          (mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_readdata),                     //                                                                   .readdata
		.F2H_Mem_Window_00000000_windowed_slave_writedata                         (mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_writedata),                    //                                                                   .writedata
		.F2H_Mem_Window_00000000_windowed_slave_burstcount                        (mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_burstcount),                   //                                                                   .burstcount
		.F2H_Mem_Window_00000000_windowed_slave_byteenable                        (mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_byteenable),                   //                                                                   .byteenable
		.F2H_Mem_Window_00000000_windowed_slave_readdatavalid                     (mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_readdatavalid),                //                                                                   .readdatavalid
		.F2H_Mem_Window_00000000_windowed_slave_waitrequest                       (mm_interconnect_0_f2h_mem_window_00000000_windowed_slave_waitrequest),                  //                                                                   .waitrequest
		.F2H_Mem_Window_FF600000_windowed_slave_address                           (mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_address),                      //                             F2H_Mem_Window_FF600000_windowed_slave.address
		.F2H_Mem_Window_FF600000_windowed_slave_write                             (mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_write),                        //                                                                   .write
		.F2H_Mem_Window_FF600000_windowed_slave_read                              (mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_read),                         //                                                                   .read
		.F2H_Mem_Window_FF600000_windowed_slave_readdata                          (mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_readdata),                     //                                                                   .readdata
		.F2H_Mem_Window_FF600000_windowed_slave_writedata                         (mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_writedata),                    //                                                                   .writedata
		.F2H_Mem_Window_FF600000_windowed_slave_burstcount                        (mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_burstcount),                   //                                                                   .burstcount
		.F2H_Mem_Window_FF600000_windowed_slave_byteenable                        (mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_byteenable),                   //                                                                   .byteenable
		.F2H_Mem_Window_FF600000_windowed_slave_readdatavalid                     (mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_readdatavalid),                //                                                                   .readdatavalid
		.F2H_Mem_Window_FF600000_windowed_slave_waitrequest                       (mm_interconnect_0_f2h_mem_window_ff600000_windowed_slave_waitrequest),                  //                                                                   .waitrequest
		.F2H_Mem_Window_FF800000_windowed_slave_address                           (mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_address),                      //                             F2H_Mem_Window_FF800000_windowed_slave.address
		.F2H_Mem_Window_FF800000_windowed_slave_write                             (mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_write),                        //                                                                   .write
		.F2H_Mem_Window_FF800000_windowed_slave_read                              (mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_read),                         //                                                                   .read
		.F2H_Mem_Window_FF800000_windowed_slave_readdata                          (mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_readdata),                     //                                                                   .readdata
		.F2H_Mem_Window_FF800000_windowed_slave_writedata                         (mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_writedata),                    //                                                                   .writedata
		.F2H_Mem_Window_FF800000_windowed_slave_burstcount                        (mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_burstcount),                   //                                                                   .burstcount
		.F2H_Mem_Window_FF800000_windowed_slave_byteenable                        (mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_byteenable),                   //                                                                   .byteenable
		.F2H_Mem_Window_FF800000_windowed_slave_readdatavalid                     (mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_readdatavalid),                //                                                                   .readdatavalid
		.F2H_Mem_Window_FF800000_windowed_slave_waitrequest                       (mm_interconnect_0_f2h_mem_window_ff800000_windowed_slave_waitrequest),                  //                                                                   .waitrequest
		.HEX3_HEX0_s1_address                                                     (mm_interconnect_0_hex3_hex0_s1_address),                                                //                                                       HEX3_HEX0_s1.address
		.HEX3_HEX0_s1_write                                                       (mm_interconnect_0_hex3_hex0_s1_write),                                                  //                                                                   .write
		.HEX3_HEX0_s1_readdata                                                    (mm_interconnect_0_hex3_hex0_s1_readdata),                                               //                                                                   .readdata
		.HEX3_HEX0_s1_writedata                                                   (mm_interconnect_0_hex3_hex0_s1_writedata),                                              //                                                                   .writedata
		.HEX3_HEX0_s1_chipselect                                                  (mm_interconnect_0_hex3_hex0_s1_chipselect),                                             //                                                                   .chipselect
		.HEX5_HEX4_s1_address                                                     (mm_interconnect_0_hex5_hex4_s1_address),                                                //                                                       HEX5_HEX4_s1.address
		.HEX5_HEX4_s1_write                                                       (mm_interconnect_0_hex5_hex4_s1_write),                                                  //                                                                   .write
		.HEX5_HEX4_s1_readdata                                                    (mm_interconnect_0_hex5_hex4_s1_readdata),                                               //                                                                   .readdata
		.HEX5_HEX4_s1_writedata                                                   (mm_interconnect_0_hex5_hex4_s1_writedata),                                              //                                                                   .writedata
		.HEX5_HEX4_s1_chipselect                                                  (mm_interconnect_0_hex5_hex4_s1_chipselect),                                             //                                                                   .chipselect
		.Interval_Timer_s1_address                                                (mm_interconnect_0_interval_timer_s1_address),                                           //                                                  Interval_Timer_s1.address
		.Interval_Timer_s1_write                                                  (mm_interconnect_0_interval_timer_s1_write),                                             //                                                                   .write
		.Interval_Timer_s1_readdata                                               (mm_interconnect_0_interval_timer_s1_readdata),                                          //                                                                   .readdata
		.Interval_Timer_s1_writedata                                              (mm_interconnect_0_interval_timer_s1_writedata),                                         //                                                                   .writedata
		.Interval_Timer_s1_chipselect                                             (mm_interconnect_0_interval_timer_s1_chipselect),                                        //                                                                   .chipselect
		.Interval_Timer_2_s1_address                                              (mm_interconnect_0_interval_timer_2_s1_address),                                         //                                                Interval_Timer_2_s1.address
		.Interval_Timer_2_s1_write                                                (mm_interconnect_0_interval_timer_2_s1_write),                                           //                                                                   .write
		.Interval_Timer_2_s1_readdata                                             (mm_interconnect_0_interval_timer_2_s1_readdata),                                        //                                                                   .readdata
		.Interval_Timer_2_s1_writedata                                            (mm_interconnect_0_interval_timer_2_s1_writedata),                                       //                                                                   .writedata
		.Interval_Timer_2_s1_chipselect                                           (mm_interconnect_0_interval_timer_2_s1_chipselect),                                      //                                                                   .chipselect
		.Interval_Timer_2nd_Core_s1_address                                       (mm_interconnect_0_interval_timer_2nd_core_s1_address),                                  //                                         Interval_Timer_2nd_Core_s1.address
		.Interval_Timer_2nd_Core_s1_write                                         (mm_interconnect_0_interval_timer_2nd_core_s1_write),                                    //                                                                   .write
		.Interval_Timer_2nd_Core_s1_readdata                                      (mm_interconnect_0_interval_timer_2nd_core_s1_readdata),                                 //                                                                   .readdata
		.Interval_Timer_2nd_Core_s1_writedata                                     (mm_interconnect_0_interval_timer_2nd_core_s1_writedata),                                //                                                                   .writedata
		.Interval_Timer_2nd_Core_s1_chipselect                                    (mm_interconnect_0_interval_timer_2nd_core_s1_chipselect),                               //                                                                   .chipselect
		.Interval_Timer_2nd_Core_2_s1_address                                     (mm_interconnect_0_interval_timer_2nd_core_2_s1_address),                                //                                       Interval_Timer_2nd_Core_2_s1.address
		.Interval_Timer_2nd_Core_2_s1_write                                       (mm_interconnect_0_interval_timer_2nd_core_2_s1_write),                                  //                                                                   .write
		.Interval_Timer_2nd_Core_2_s1_readdata                                    (mm_interconnect_0_interval_timer_2nd_core_2_s1_readdata),                               //                                                                   .readdata
		.Interval_Timer_2nd_Core_2_s1_writedata                                   (mm_interconnect_0_interval_timer_2nd_core_2_s1_writedata),                              //                                                                   .writedata
		.Interval_Timer_2nd_Core_2_s1_chipselect                                  (mm_interconnect_0_interval_timer_2nd_core_2_s1_chipselect),                             //                                                                   .chipselect
		.IrDA_avalon_irda_slave_address                                           (mm_interconnect_0_irda_avalon_irda_slave_address),                                      //                                             IrDA_avalon_irda_slave.address
		.IrDA_avalon_irda_slave_write                                             (mm_interconnect_0_irda_avalon_irda_slave_write),                                        //                                                                   .write
		.IrDA_avalon_irda_slave_read                                              (mm_interconnect_0_irda_avalon_irda_slave_read),                                         //                                                                   .read
		.IrDA_avalon_irda_slave_readdata                                          (mm_interconnect_0_irda_avalon_irda_slave_readdata),                                     //                                                                   .readdata
		.IrDA_avalon_irda_slave_writedata                                         (mm_interconnect_0_irda_avalon_irda_slave_writedata),                                    //                                                                   .writedata
		.IrDA_avalon_irda_slave_byteenable                                        (mm_interconnect_0_irda_avalon_irda_slave_byteenable),                                   //                                                                   .byteenable
		.IrDA_avalon_irda_slave_chipselect                                        (mm_interconnect_0_irda_avalon_irda_slave_chipselect),                                   //                                                                   .chipselect
		.JTAG_UART_avalon_jtag_slave_address                                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                                 //                                        JTAG_UART_avalon_jtag_slave.address
		.JTAG_UART_avalon_jtag_slave_write                                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                                   //                                                                   .write
		.JTAG_UART_avalon_jtag_slave_read                                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                                    //                                                                   .read
		.JTAG_UART_avalon_jtag_slave_readdata                                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),                                //                                                                   .readdata
		.JTAG_UART_avalon_jtag_slave_writedata                                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),                               //                                                                   .writedata
		.JTAG_UART_avalon_jtag_slave_waitrequest                                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),                             //                                                                   .waitrequest
		.JTAG_UART_avalon_jtag_slave_chipselect                                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),                              //                                                                   .chipselect
		.JTAG_UART_2nd_Core_avalon_jtag_slave_address                             (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_address),                        //                               JTAG_UART_2nd_Core_avalon_jtag_slave.address
		.JTAG_UART_2nd_Core_avalon_jtag_slave_write                               (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write),                          //                                                                   .write
		.JTAG_UART_2nd_Core_avalon_jtag_slave_read                                (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read),                           //                                                                   .read
		.JTAG_UART_2nd_Core_avalon_jtag_slave_readdata                            (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_readdata),                       //                                                                   .readdata
		.JTAG_UART_2nd_Core_avalon_jtag_slave_writedata                           (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_writedata),                      //                                                                   .writedata
		.JTAG_UART_2nd_Core_avalon_jtag_slave_waitrequest                         (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_waitrequest),                    //                                                                   .waitrequest
		.JTAG_UART_2nd_Core_avalon_jtag_slave_chipselect                          (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_chipselect),                     //                                                                   .chipselect
		.JTAG_UART_for_ARM_0_avalon_jtag_slave_address                            (mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_address),                       //                              JTAG_UART_for_ARM_0_avalon_jtag_slave.address
		.JTAG_UART_for_ARM_0_avalon_jtag_slave_write                              (mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_write),                         //                                                                   .write
		.JTAG_UART_for_ARM_0_avalon_jtag_slave_read                               (mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_read),                          //                                                                   .read
		.JTAG_UART_for_ARM_0_avalon_jtag_slave_readdata                           (mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_readdata),                      //                                                                   .readdata
		.JTAG_UART_for_ARM_0_avalon_jtag_slave_writedata                          (mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_writedata),                     //                                                                   .writedata
		.JTAG_UART_for_ARM_0_avalon_jtag_slave_waitrequest                        (mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_waitrequest),                   //                                                                   .waitrequest
		.JTAG_UART_for_ARM_0_avalon_jtag_slave_chipselect                         (mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_chipselect),                    //                                                                   .chipselect
		.JTAG_UART_for_ARM_1_avalon_jtag_slave_address                            (mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_address),                       //                              JTAG_UART_for_ARM_1_avalon_jtag_slave.address
		.JTAG_UART_for_ARM_1_avalon_jtag_slave_write                              (mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_write),                         //                                                                   .write
		.JTAG_UART_for_ARM_1_avalon_jtag_slave_read                               (mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_read),                          //                                                                   .read
		.JTAG_UART_for_ARM_1_avalon_jtag_slave_readdata                           (mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_readdata),                      //                                                                   .readdata
		.JTAG_UART_for_ARM_1_avalon_jtag_slave_writedata                          (mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_writedata),                     //                                                                   .writedata
		.JTAG_UART_for_ARM_1_avalon_jtag_slave_waitrequest                        (mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_waitrequest),                   //                                                                   .waitrequest
		.JTAG_UART_for_ARM_1_avalon_jtag_slave_chipselect                         (mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_chipselect),                    //                                                                   .chipselect
		.LEDs_s1_address                                                          (mm_interconnect_0_leds_s1_address),                                                     //                                                            LEDs_s1.address
		.LEDs_s1_write                                                            (mm_interconnect_0_leds_s1_write),                                                       //                                                                   .write
		.LEDs_s1_readdata                                                         (mm_interconnect_0_leds_s1_readdata),                                                    //                                                                   .readdata
		.LEDs_s1_writedata                                                        (mm_interconnect_0_leds_s1_writedata),                                                   //                                                                   .writedata
		.LEDs_s1_chipselect                                                       (mm_interconnect_0_leds_s1_chipselect),                                                  //                                                                   .chipselect
		.Nios2_debug_mem_slave_address                                            (mm_interconnect_0_nios2_debug_mem_slave_address),                                       //                                              Nios2_debug_mem_slave.address
		.Nios2_debug_mem_slave_write                                              (mm_interconnect_0_nios2_debug_mem_slave_write),                                         //                                                                   .write
		.Nios2_debug_mem_slave_read                                               (mm_interconnect_0_nios2_debug_mem_slave_read),                                          //                                                                   .read
		.Nios2_debug_mem_slave_readdata                                           (mm_interconnect_0_nios2_debug_mem_slave_readdata),                                      //                                                                   .readdata
		.Nios2_debug_mem_slave_writedata                                          (mm_interconnect_0_nios2_debug_mem_slave_writedata),                                     //                                                                   .writedata
		.Nios2_debug_mem_slave_byteenable                                         (mm_interconnect_0_nios2_debug_mem_slave_byteenable),                                    //                                                                   .byteenable
		.Nios2_debug_mem_slave_waitrequest                                        (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),                                   //                                                                   .waitrequest
		.Nios2_debug_mem_slave_debugaccess                                        (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),                                   //                                                                   .debugaccess
		.Nios2_2nd_Core_debug_mem_slave_address                                   (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_address),                              //                                     Nios2_2nd_Core_debug_mem_slave.address
		.Nios2_2nd_Core_debug_mem_slave_write                                     (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_write),                                //                                                                   .write
		.Nios2_2nd_Core_debug_mem_slave_read                                      (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_read),                                 //                                                                   .read
		.Nios2_2nd_Core_debug_mem_slave_readdata                                  (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_readdata),                             //                                                                   .readdata
		.Nios2_2nd_Core_debug_mem_slave_writedata                                 (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_writedata),                            //                                                                   .writedata
		.Nios2_2nd_Core_debug_mem_slave_byteenable                                (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_byteenable),                           //                                                                   .byteenable
		.Nios2_2nd_Core_debug_mem_slave_waitrequest                               (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_waitrequest),                          //                                                                   .waitrequest
		.Nios2_2nd_Core_debug_mem_slave_debugaccess                               (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_debugaccess),                          //                                                                   .debugaccess
		.Onchip_SRAM_s1_address                                                   (mm_interconnect_0_onchip_sram_s1_address),                                              //                                                     Onchip_SRAM_s1.address
		.Onchip_SRAM_s1_write                                                     (mm_interconnect_0_onchip_sram_s1_write),                                                //                                                                   .write
		.Onchip_SRAM_s1_readdata                                                  (mm_interconnect_0_onchip_sram_s1_readdata),                                             //                                                                   .readdata
		.Onchip_SRAM_s1_writedata                                                 (mm_interconnect_0_onchip_sram_s1_writedata),                                            //                                                                   .writedata
		.Onchip_SRAM_s1_byteenable                                                (mm_interconnect_0_onchip_sram_s1_byteenable),                                           //                                                                   .byteenable
		.Onchip_SRAM_s1_chipselect                                                (mm_interconnect_0_onchip_sram_s1_chipselect),                                           //                                                                   .chipselect
		.Onchip_SRAM_s1_clken                                                     (mm_interconnect_0_onchip_sram_s1_clken),                                                //                                                                   .clken
		.Onchip_SRAM_s2_address                                                   (mm_interconnect_0_onchip_sram_s2_address),                                              //                                                     Onchip_SRAM_s2.address
		.Onchip_SRAM_s2_write                                                     (mm_interconnect_0_onchip_sram_s2_write),                                                //                                                                   .write
		.Onchip_SRAM_s2_readdata                                                  (mm_interconnect_0_onchip_sram_s2_readdata),                                             //                                                                   .readdata
		.Onchip_SRAM_s2_writedata                                                 (mm_interconnect_0_onchip_sram_s2_writedata),                                            //                                                                   .writedata
		.Onchip_SRAM_s2_byteenable                                                (mm_interconnect_0_onchip_sram_s2_byteenable),                                           //                                                                   .byteenable
		.Onchip_SRAM_s2_chipselect                                                (mm_interconnect_0_onchip_sram_s2_chipselect),                                           //                                                                   .chipselect
		.Onchip_SRAM_s2_clken                                                     (mm_interconnect_0_onchip_sram_s2_clken),                                                //                                                                   .clken
		.Pixel_DMA_Addr_Translation_slave_address                                 (mm_interconnect_0_pixel_dma_addr_translation_slave_address),                            //                                   Pixel_DMA_Addr_Translation_slave.address
		.Pixel_DMA_Addr_Translation_slave_write                                   (mm_interconnect_0_pixel_dma_addr_translation_slave_write),                              //                                                                   .write
		.Pixel_DMA_Addr_Translation_slave_read                                    (mm_interconnect_0_pixel_dma_addr_translation_slave_read),                               //                                                                   .read
		.Pixel_DMA_Addr_Translation_slave_readdata                                (mm_interconnect_0_pixel_dma_addr_translation_slave_readdata),                           //                                                                   .readdata
		.Pixel_DMA_Addr_Translation_slave_writedata                               (mm_interconnect_0_pixel_dma_addr_translation_slave_writedata),                          //                                                                   .writedata
		.Pixel_DMA_Addr_Translation_slave_byteenable                              (mm_interconnect_0_pixel_dma_addr_translation_slave_byteenable),                         //                                                                   .byteenable
		.Pixel_DMA_Addr_Translation_slave_waitrequest                             (mm_interconnect_0_pixel_dma_addr_translation_slave_waitrequest),                        //                                                                   .waitrequest
		.PS2_Port_avalon_ps2_slave_address                                        (mm_interconnect_0_ps2_port_avalon_ps2_slave_address),                                   //                                          PS2_Port_avalon_ps2_slave.address
		.PS2_Port_avalon_ps2_slave_write                                          (mm_interconnect_0_ps2_port_avalon_ps2_slave_write),                                     //                                                                   .write
		.PS2_Port_avalon_ps2_slave_read                                           (mm_interconnect_0_ps2_port_avalon_ps2_slave_read),                                      //                                                                   .read
		.PS2_Port_avalon_ps2_slave_readdata                                       (mm_interconnect_0_ps2_port_avalon_ps2_slave_readdata),                                  //                                                                   .readdata
		.PS2_Port_avalon_ps2_slave_writedata                                      (mm_interconnect_0_ps2_port_avalon_ps2_slave_writedata),                                 //                                                                   .writedata
		.PS2_Port_avalon_ps2_slave_byteenable                                     (mm_interconnect_0_ps2_port_avalon_ps2_slave_byteenable),                                //                                                                   .byteenable
		.PS2_Port_avalon_ps2_slave_waitrequest                                    (mm_interconnect_0_ps2_port_avalon_ps2_slave_waitrequest),                               //                                                                   .waitrequest
		.PS2_Port_avalon_ps2_slave_chipselect                                     (mm_interconnect_0_ps2_port_avalon_ps2_slave_chipselect),                                //                                                                   .chipselect
		.PS2_Port_Dual_avalon_ps2_slave_address                                   (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_address),                              //                                     PS2_Port_Dual_avalon_ps2_slave.address
		.PS2_Port_Dual_avalon_ps2_slave_write                                     (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_write),                                //                                                                   .write
		.PS2_Port_Dual_avalon_ps2_slave_read                                      (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_read),                                 //                                                                   .read
		.PS2_Port_Dual_avalon_ps2_slave_readdata                                  (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_readdata),                             //                                                                   .readdata
		.PS2_Port_Dual_avalon_ps2_slave_writedata                                 (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_writedata),                            //                                                                   .writedata
		.PS2_Port_Dual_avalon_ps2_slave_byteenable                                (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_byteenable),                           //                                                                   .byteenable
		.PS2_Port_Dual_avalon_ps2_slave_waitrequest                               (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_waitrequest),                          //                                                                   .waitrequest
		.PS2_Port_Dual_avalon_ps2_slave_chipselect                                (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_chipselect),                           //                                                                   .chipselect
		.Pushbuttons_s1_address                                                   (mm_interconnect_0_pushbuttons_s1_address),                                              //                                                     Pushbuttons_s1.address
		.Pushbuttons_s1_write                                                     (mm_interconnect_0_pushbuttons_s1_write),                                                //                                                                   .write
		.Pushbuttons_s1_readdata                                                  (mm_interconnect_0_pushbuttons_s1_readdata),                                             //                                                                   .readdata
		.Pushbuttons_s1_writedata                                                 (mm_interconnect_0_pushbuttons_s1_writedata),                                            //                                                                   .writedata
		.Pushbuttons_s1_chipselect                                                (mm_interconnect_0_pushbuttons_s1_chipselect),                                           //                                                                   .chipselect
		.SDRAM_s1_address                                                         (mm_interconnect_0_sdram_s1_address),                                                    //                                                           SDRAM_s1.address
		.SDRAM_s1_write                                                           (mm_interconnect_0_sdram_s1_write),                                                      //                                                                   .write
		.SDRAM_s1_read                                                            (mm_interconnect_0_sdram_s1_read),                                                       //                                                                   .read
		.SDRAM_s1_readdata                                                        (mm_interconnect_0_sdram_s1_readdata),                                                   //                                                                   .readdata
		.SDRAM_s1_writedata                                                       (mm_interconnect_0_sdram_s1_writedata),                                                  //                                                                   .writedata
		.SDRAM_s1_byteenable                                                      (mm_interconnect_0_sdram_s1_byteenable),                                                 //                                                                   .byteenable
		.SDRAM_s1_readdatavalid                                                   (mm_interconnect_0_sdram_s1_readdatavalid),                                              //                                                                   .readdatavalid
		.SDRAM_s1_waitrequest                                                     (mm_interconnect_0_sdram_s1_waitrequest),                                                //                                                                   .waitrequest
		.SDRAM_s1_chipselect                                                      (mm_interconnect_0_sdram_s1_chipselect),                                                 //                                                                   .chipselect
		.Slider_Switches_s1_address                                               (mm_interconnect_0_slider_switches_s1_address),                                          //                                                 Slider_Switches_s1.address
		.Slider_Switches_s1_readdata                                              (mm_interconnect_0_slider_switches_s1_readdata),                                         //                                                                   .readdata
		.SysID_control_slave_address                                              (mm_interconnect_0_sysid_control_slave_address),                                         //                                                SysID_control_slave.address
		.SysID_control_slave_readdata                                             (mm_interconnect_0_sysid_control_slave_readdata),                                        //                                                                   .readdata
		.VGA_Subsystem_char_buffer_control_slave_address                          (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_address),                     //                            VGA_Subsystem_char_buffer_control_slave.address
		.VGA_Subsystem_char_buffer_control_slave_write                            (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_write),                       //                                                                   .write
		.VGA_Subsystem_char_buffer_control_slave_read                             (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_read),                        //                                                                   .read
		.VGA_Subsystem_char_buffer_control_slave_readdata                         (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_readdata),                    //                                                                   .readdata
		.VGA_Subsystem_char_buffer_control_slave_writedata                        (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_writedata),                   //                                                                   .writedata
		.VGA_Subsystem_char_buffer_control_slave_byteenable                       (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_byteenable),                  //                                                                   .byteenable
		.VGA_Subsystem_char_buffer_slave_address                                  (mm_interconnect_0_vga_subsystem_char_buffer_slave_address),                             //                                    VGA_Subsystem_char_buffer_slave.address
		.VGA_Subsystem_char_buffer_slave_write                                    (mm_interconnect_0_vga_subsystem_char_buffer_slave_write),                               //                                                                   .write
		.VGA_Subsystem_char_buffer_slave_readdata                                 (mm_interconnect_0_vga_subsystem_char_buffer_slave_readdata),                            //                                                                   .readdata
		.VGA_Subsystem_char_buffer_slave_writedata                                (mm_interconnect_0_vga_subsystem_char_buffer_slave_writedata),                           //                                                                   .writedata
		.VGA_Subsystem_char_buffer_slave_byteenable                               (mm_interconnect_0_vga_subsystem_char_buffer_slave_byteenable),                          //                                                                   .byteenable
		.VGA_Subsystem_char_buffer_slave_chipselect                               (mm_interconnect_0_vga_subsystem_char_buffer_slave_chipselect),                          //                                                                   .chipselect
		.VGA_Subsystem_char_buffer_slave_clken                                    (mm_interconnect_0_vga_subsystem_char_buffer_slave_clken),                               //                                                                   .clken
		.VGA_Subsystem_pixel_dma_control_slave_address                            (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_address),                       //                              VGA_Subsystem_pixel_dma_control_slave.address
		.VGA_Subsystem_pixel_dma_control_slave_write                              (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_write),                         //                                                                   .write
		.VGA_Subsystem_pixel_dma_control_slave_read                               (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_read),                          //                                                                   .read
		.VGA_Subsystem_pixel_dma_control_slave_readdata                           (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_readdata),                      //                                                                   .readdata
		.VGA_Subsystem_pixel_dma_control_slave_writedata                          (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_writedata),                     //                                                                   .writedata
		.VGA_Subsystem_pixel_dma_control_slave_byteenable                         (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_byteenable),                    //                                                                   .byteenable
		.VGA_Subsystem_rgb_slave_read                                             (mm_interconnect_0_vga_subsystem_rgb_slave_read),                                        //                                            VGA_Subsystem_rgb_slave.read
		.VGA_Subsystem_rgb_slave_readdata                                         (mm_interconnect_0_vga_subsystem_rgb_slave_readdata),                                    //                                                                   .readdata
		.Video_In_DMA_Addr_Translation_slave_address                              (mm_interconnect_0_video_in_dma_addr_translation_slave_address),                         //                                Video_In_DMA_Addr_Translation_slave.address
		.Video_In_DMA_Addr_Translation_slave_write                                (mm_interconnect_0_video_in_dma_addr_translation_slave_write),                           //                                                                   .write
		.Video_In_DMA_Addr_Translation_slave_read                                 (mm_interconnect_0_video_in_dma_addr_translation_slave_read),                            //                                                                   .read
		.Video_In_DMA_Addr_Translation_slave_readdata                             (mm_interconnect_0_video_in_dma_addr_translation_slave_readdata),                        //                                                                   .readdata
		.Video_In_DMA_Addr_Translation_slave_writedata                            (mm_interconnect_0_video_in_dma_addr_translation_slave_writedata),                       //                                                                   .writedata
		.Video_In_DMA_Addr_Translation_slave_byteenable                           (mm_interconnect_0_video_in_dma_addr_translation_slave_byteenable),                      //                                                                   .byteenable
		.Video_In_DMA_Addr_Translation_slave_waitrequest                          (mm_interconnect_0_video_in_dma_addr_translation_slave_waitrequest),                     //                                                                   .waitrequest
		.Video_In_Subsystem_video_in_dma_control_slave_address                    (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_address),               //                      Video_In_Subsystem_video_in_dma_control_slave.address
		.Video_In_Subsystem_video_in_dma_control_slave_write                      (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_write),                 //                                                                   .write
		.Video_In_Subsystem_video_in_dma_control_slave_read                       (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_read),                  //                                                                   .read
		.Video_In_Subsystem_video_in_dma_control_slave_readdata                   (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_readdata),              //                                                                   .readdata
		.Video_In_Subsystem_video_in_dma_control_slave_writedata                  (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_writedata),             //                                                                   .writedata
		.Video_In_Subsystem_video_in_dma_control_slave_byteenable                 (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_byteenable),            //                                                                   .byteenable
		.Video_In_Subsystem_video_in_edge_detection_control_slave_address         (mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_address),    //           Video_In_Subsystem_video_in_edge_detection_control_slave.address
		.Video_In_Subsystem_video_in_edge_detection_control_slave_write           (mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_write),      //                                                                   .write
		.Video_In_Subsystem_video_in_edge_detection_control_slave_readdata        (mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_readdata),   //                                                                   .readdata
		.Video_In_Subsystem_video_in_edge_detection_control_slave_writedata       (mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_writedata),  //                                                                   .writedata
		.Video_In_Subsystem_video_in_edge_detection_control_slave_chipselect      (mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_chipselect)  //                                                                   .chipselect
	);

	Computer_System_mm_interconnect_1 mm_interconnect_1 (
		.ARM_A9_HPS_f2h_axi_slave_awid                                         (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awid),       //                                        ARM_A9_HPS_f2h_axi_slave.awid
		.ARM_A9_HPS_f2h_axi_slave_awaddr                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awaddr),     //                                                                .awaddr
		.ARM_A9_HPS_f2h_axi_slave_awlen                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlen),      //                                                                .awlen
		.ARM_A9_HPS_f2h_axi_slave_awsize                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awsize),     //                                                                .awsize
		.ARM_A9_HPS_f2h_axi_slave_awburst                                      (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awburst),    //                                                                .awburst
		.ARM_A9_HPS_f2h_axi_slave_awlock                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlock),     //                                                                .awlock
		.ARM_A9_HPS_f2h_axi_slave_awcache                                      (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awcache),    //                                                                .awcache
		.ARM_A9_HPS_f2h_axi_slave_awprot                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awprot),     //                                                                .awprot
		.ARM_A9_HPS_f2h_axi_slave_awuser                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awuser),     //                                                                .awuser
		.ARM_A9_HPS_f2h_axi_slave_awvalid                                      (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awvalid),    //                                                                .awvalid
		.ARM_A9_HPS_f2h_axi_slave_awready                                      (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awready),    //                                                                .awready
		.ARM_A9_HPS_f2h_axi_slave_wid                                          (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wid),        //                                                                .wid
		.ARM_A9_HPS_f2h_axi_slave_wdata                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wdata),      //                                                                .wdata
		.ARM_A9_HPS_f2h_axi_slave_wstrb                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wstrb),      //                                                                .wstrb
		.ARM_A9_HPS_f2h_axi_slave_wlast                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wlast),      //                                                                .wlast
		.ARM_A9_HPS_f2h_axi_slave_wvalid                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wvalid),     //                                                                .wvalid
		.ARM_A9_HPS_f2h_axi_slave_wready                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wready),     //                                                                .wready
		.ARM_A9_HPS_f2h_axi_slave_bid                                          (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bid),        //                                                                .bid
		.ARM_A9_HPS_f2h_axi_slave_bresp                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bresp),      //                                                                .bresp
		.ARM_A9_HPS_f2h_axi_slave_bvalid                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bvalid),     //                                                                .bvalid
		.ARM_A9_HPS_f2h_axi_slave_bready                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bready),     //                                                                .bready
		.ARM_A9_HPS_f2h_axi_slave_arid                                         (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arid),       //                                                                .arid
		.ARM_A9_HPS_f2h_axi_slave_araddr                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_araddr),     //                                                                .araddr
		.ARM_A9_HPS_f2h_axi_slave_arlen                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlen),      //                                                                .arlen
		.ARM_A9_HPS_f2h_axi_slave_arsize                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arsize),     //                                                                .arsize
		.ARM_A9_HPS_f2h_axi_slave_arburst                                      (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arburst),    //                                                                .arburst
		.ARM_A9_HPS_f2h_axi_slave_arlock                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlock),     //                                                                .arlock
		.ARM_A9_HPS_f2h_axi_slave_arcache                                      (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arcache),    //                                                                .arcache
		.ARM_A9_HPS_f2h_axi_slave_arprot                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arprot),     //                                                                .arprot
		.ARM_A9_HPS_f2h_axi_slave_aruser                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_aruser),     //                                                                .aruser
		.ARM_A9_HPS_f2h_axi_slave_arvalid                                      (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arvalid),    //                                                                .arvalid
		.ARM_A9_HPS_f2h_axi_slave_arready                                      (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arready),    //                                                                .arready
		.ARM_A9_HPS_f2h_axi_slave_rid                                          (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rid),        //                                                                .rid
		.ARM_A9_HPS_f2h_axi_slave_rdata                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rdata),      //                                                                .rdata
		.ARM_A9_HPS_f2h_axi_slave_rresp                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rresp),      //                                                                .rresp
		.ARM_A9_HPS_f2h_axi_slave_rlast                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rlast),      //                                                                .rlast
		.ARM_A9_HPS_f2h_axi_slave_rvalid                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rvalid),     //                                                                .rvalid
		.ARM_A9_HPS_f2h_axi_slave_rready                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rready),     //                                                                .rready
		.System_PLL_sys_clk_clk                                                (system_pll_sys_clk_clk),                                //                                              System_PLL_sys_clk.clk
		.ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset (rst_controller_008_reset_out_reset),                    // ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.F2H_Mem_Window_00000000_reset_reset_bridge_in_reset_reset             (rst_controller_reset_out_reset),                        //             F2H_Mem_Window_00000000_reset_reset_bridge_in_reset.reset
		.JTAG_to_HPS_Bridge_clk_reset_reset_bridge_in_reset_reset              (rst_controller_reset_out_reset),                        //              JTAG_to_HPS_Bridge_clk_reset_reset_bridge_in_reset.reset
		.F2H_Mem_Window_00000000_expanded_master_address                       (f2h_mem_window_00000000_expanded_master_address),       //                         F2H_Mem_Window_00000000_expanded_master.address
		.F2H_Mem_Window_00000000_expanded_master_waitrequest                   (f2h_mem_window_00000000_expanded_master_waitrequest),   //                                                                .waitrequest
		.F2H_Mem_Window_00000000_expanded_master_burstcount                    (f2h_mem_window_00000000_expanded_master_burstcount),    //                                                                .burstcount
		.F2H_Mem_Window_00000000_expanded_master_byteenable                    (f2h_mem_window_00000000_expanded_master_byteenable),    //                                                                .byteenable
		.F2H_Mem_Window_00000000_expanded_master_read                          (f2h_mem_window_00000000_expanded_master_read),          //                                                                .read
		.F2H_Mem_Window_00000000_expanded_master_readdata                      (f2h_mem_window_00000000_expanded_master_readdata),      //                                                                .readdata
		.F2H_Mem_Window_00000000_expanded_master_readdatavalid                 (f2h_mem_window_00000000_expanded_master_readdatavalid), //                                                                .readdatavalid
		.F2H_Mem_Window_00000000_expanded_master_write                         (f2h_mem_window_00000000_expanded_master_write),         //                                                                .write
		.F2H_Mem_Window_00000000_expanded_master_writedata                     (f2h_mem_window_00000000_expanded_master_writedata),     //                                                                .writedata
		.F2H_Mem_Window_FF600000_expanded_master_address                       (f2h_mem_window_ff600000_expanded_master_address),       //                         F2H_Mem_Window_FF600000_expanded_master.address
		.F2H_Mem_Window_FF600000_expanded_master_waitrequest                   (f2h_mem_window_ff600000_expanded_master_waitrequest),   //                                                                .waitrequest
		.F2H_Mem_Window_FF600000_expanded_master_burstcount                    (f2h_mem_window_ff600000_expanded_master_burstcount),    //                                                                .burstcount
		.F2H_Mem_Window_FF600000_expanded_master_byteenable                    (f2h_mem_window_ff600000_expanded_master_byteenable),    //                                                                .byteenable
		.F2H_Mem_Window_FF600000_expanded_master_read                          (f2h_mem_window_ff600000_expanded_master_read),          //                                                                .read
		.F2H_Mem_Window_FF600000_expanded_master_readdata                      (f2h_mem_window_ff600000_expanded_master_readdata),      //                                                                .readdata
		.F2H_Mem_Window_FF600000_expanded_master_readdatavalid                 (f2h_mem_window_ff600000_expanded_master_readdatavalid), //                                                                .readdatavalid
		.F2H_Mem_Window_FF600000_expanded_master_write                         (f2h_mem_window_ff600000_expanded_master_write),         //                                                                .write
		.F2H_Mem_Window_FF600000_expanded_master_writedata                     (f2h_mem_window_ff600000_expanded_master_writedata),     //                                                                .writedata
		.F2H_Mem_Window_FF800000_expanded_master_address                       (f2h_mem_window_ff800000_expanded_master_address),       //                         F2H_Mem_Window_FF800000_expanded_master.address
		.F2H_Mem_Window_FF800000_expanded_master_waitrequest                   (f2h_mem_window_ff800000_expanded_master_waitrequest),   //                                                                .waitrequest
		.F2H_Mem_Window_FF800000_expanded_master_burstcount                    (f2h_mem_window_ff800000_expanded_master_burstcount),    //                                                                .burstcount
		.F2H_Mem_Window_FF800000_expanded_master_byteenable                    (f2h_mem_window_ff800000_expanded_master_byteenable),    //                                                                .byteenable
		.F2H_Mem_Window_FF800000_expanded_master_read                          (f2h_mem_window_ff800000_expanded_master_read),          //                                                                .read
		.F2H_Mem_Window_FF800000_expanded_master_readdata                      (f2h_mem_window_ff800000_expanded_master_readdata),      //                                                                .readdata
		.F2H_Mem_Window_FF800000_expanded_master_readdatavalid                 (f2h_mem_window_ff800000_expanded_master_readdatavalid), //                                                                .readdatavalid
		.F2H_Mem_Window_FF800000_expanded_master_write                         (f2h_mem_window_ff800000_expanded_master_write),         //                                                                .write
		.F2H_Mem_Window_FF800000_expanded_master_writedata                     (f2h_mem_window_ff800000_expanded_master_writedata),     //                                                                .writedata
		.JTAG_to_HPS_Bridge_master_address                                     (jtag_to_hps_bridge_master_address),                     //                                       JTAG_to_HPS_Bridge_master.address
		.JTAG_to_HPS_Bridge_master_waitrequest                                 (jtag_to_hps_bridge_master_waitrequest),                 //                                                                .waitrequest
		.JTAG_to_HPS_Bridge_master_byteenable                                  (jtag_to_hps_bridge_master_byteenable),                  //                                                                .byteenable
		.JTAG_to_HPS_Bridge_master_read                                        (jtag_to_hps_bridge_master_read),                        //                                                                .read
		.JTAG_to_HPS_Bridge_master_readdata                                    (jtag_to_hps_bridge_master_readdata),                    //                                                                .readdata
		.JTAG_to_HPS_Bridge_master_readdatavalid                               (jtag_to_hps_bridge_master_readdatavalid),               //                                                                .readdatavalid
		.JTAG_to_HPS_Bridge_master_write                                       (jtag_to_hps_bridge_master_write),                       //                                                                .write
		.JTAG_to_HPS_Bridge_master_writedata                                   (jtag_to_hps_bridge_master_writedata)                    //                                                                .writedata
	);

	Computer_System_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq), // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq), // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq), // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq), // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq), // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq), // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq), // receiver7.irq
		.receiver8_irq (irq_mapper_receiver8_irq), // receiver8.irq
		.sender_irq    (arm_a9_hps_f2h_irq0_irq)   //    sender.irq
	);

	Computer_System_irq_mapper_001 irq_mapper_001 (
		.clk           (),                             //       clk.clk
		.reset         (),                             // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq), // receiver0.irq
		.sender_irq    (arm_a9_hps_f2h_irq1_irq)       //    sender.irq
	);

	Computer_System_irq_mapper irq_mapper_002 (
		.clk           (system_pll_sys_clk_clk),             //       clk.clk
		.reset         (rst_controller_004_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.receiver6_irq (irq_mapper_002_receiver6_irq),       // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),           // receiver7.irq
		.receiver8_irq (irq_mapper_receiver8_irq),           // receiver8.irq
		.sender_irq    (nios2_irq_irq)                       //    sender.irq
	);

	Computer_System_irq_mapper irq_mapper_003 (
		.clk           (system_pll_sys_clk_clk),             //       clk.clk
		.reset         (rst_controller_005_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.receiver6_irq (irq_mapper_003_receiver6_irq),       // receiver6.irq
		.receiver7_irq (irq_mapper_003_receiver7_irq),       // receiver7.irq
		.receiver8_irq (irq_mapper_003_receiver8_irq),       // receiver8.irq
		.sender_irq    (nios2_2nd_core_irq_irq)              //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (nios2_debug_reset_request_reset),    // reset_in0.reset
		.reset_in1      (~arm_a9_hps_h2f_reset_reset),        // reset_in1.reset
		.reset_in2      (system_pll_reset_source_reset),      // reset_in2.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (nios2_2nd_core_debug_reset_request_reset), // reset_in0.reset
		.reset_in1      (~arm_a9_hps_h2f_reset_reset),              // reset_in1.reset
		.reset_in2      (system_pll_reset_source_reset),            // reset_in2.reset
		.clk            (system_pll_sys_clk_clk),                   //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset),       // reset_out.reset
		.reset_req      (),                                         // (terminated)
		.reset_req_in0  (1'b0),                                     // (terminated)
		.reset_req_in1  (1'b0),                                     // (terminated)
		.reset_req_in2  (1'b0),                                     // (terminated)
		.reset_in3      (1'b0),                                     // (terminated)
		.reset_req_in3  (1'b0),                                     // (terminated)
		.reset_in4      (1'b0),                                     // (terminated)
		.reset_req_in4  (1'b0),                                     // (terminated)
		.reset_in5      (1'b0),                                     // (terminated)
		.reset_req_in5  (1'b0),                                     // (terminated)
		.reset_in6      (1'b0),                                     // (terminated)
		.reset_req_in6  (1'b0),                                     // (terminated)
		.reset_in7      (1'b0),                                     // (terminated)
		.reset_req_in7  (1'b0),                                     // (terminated)
		.reset_in8      (1'b0),                                     // (terminated)
		.reset_req_in8  (1'b0),                                     // (terminated)
		.reset_in9      (1'b0),                                     // (terminated)
		.reset_req_in9  (1'b0),                                     // (terminated)
		.reset_in10     (1'b0),                                     // (terminated)
		.reset_req_in10 (1'b0),                                     // (terminated)
		.reset_in11     (1'b0),                                     // (terminated)
		.reset_req_in11 (1'b0),                                     // (terminated)
		.reset_in12     (1'b0),                                     // (terminated)
		.reset_req_in12 (1'b0),                                     // (terminated)
		.reset_in13     (1'b0),                                     // (terminated)
		.reset_req_in13 (1'b0),                                     // (terminated)
		.reset_in14     (1'b0),                                     // (terminated)
		.reset_req_in14 (1'b0),                                     // (terminated)
		.reset_in15     (1'b0),                                     // (terminated)
		.reset_req_in15 (1'b0)                                      // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_007 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_007_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_008 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_008_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
